module front_panel_interface
(
	input wire clk, reset,
	input wire[9:0] disp_w,	         // Display brightness
	input wire disp_en,              // Display enable
	
	
	
);

endmodule