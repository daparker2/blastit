// controller_tb.v

// Generated using ACDS version 13.1 162 at 2018.07.11.00:25:35

`timescale 1 ps / 1 ps
module controller_tb (
	);

	wire         controller_inst_clk_bfm_clk_clk;                   // controller_inst_clk_bfm:clk -> controller_inst:clk_clk
	wire   [7:0] controller_inst_command_tx_export;                 // controller_inst:command_tx_export -> controller_inst_command_tx_bfm:sig_export
	wire   [7:0] controller_inst_command_rx_bfm_conduit_export;     // controller_inst_command_rx_bfm:sig_export -> controller_inst:command_rx_export
	wire   [7:0] controller_inst_command_status_bfm_conduit_export; // controller_inst_command_status_bfm:sig_export -> controller_inst:command_status_export
	wire   [8:0] controller_inst_disp_en_brightness_export;         // controller_inst:disp_en_brightness_export -> controller_inst_disp_en_brightness_bfm:sig_export
	wire   [2:0] controller_inst_system_status_bfm_conduit_export;  // controller_inst_system_status_bfm:sig_export -> controller_inst:system_status_export
	wire   [1:0] controller_inst_command_en_export;                 // controller_inst:command_en_export -> controller_inst_command_en_bfm:sig_export
	wire   [2:0] controller_inst_warning_en_export;                 // controller_inst:warning_en_export -> controller_inst_warning_en_bfm:sig_export
	wire  [11:0] controller_inst_boost_export;                      // controller_inst:boost_export -> controller_inst_boost_bfm:sig_export
	wire  [11:0] controller_inst_afr_export;                        // controller_inst:afr_export -> controller_inst_afr_bfm:sig_export
	wire  [11:0] controller_inst_oil_temp_export;                   // controller_inst:oil_temp_export -> controller_inst_oil_temp_bfm:sig_export
	wire  [11:0] controller_inst_coolant_temp_export;               // controller_inst:coolant_temp_export -> controller_inst_coolant_temp_bfm:sig_export
	wire  [11:0] controller_inst_intake_temp_export;                // controller_inst:intake_temp_export -> controller_inst_intake_temp_bfm:sig_export
	wire         controller_inst_ign_en_export;                     // controller_inst:ign_en_export -> controller_inst_ign_en_bfm:sig_export

	controller controller_inst (
		.clk_clk                   (controller_inst_clk_bfm_clk_clk),                   //                clk.clk
		.command_tx_export         (controller_inst_command_tx_export),                 //         command_tx.export
		.command_rx_export         (controller_inst_command_rx_bfm_conduit_export),     //         command_rx.export
		.command_status_export     (controller_inst_command_status_bfm_conduit_export), //     command_status.export
		.disp_en_brightness_export (controller_inst_disp_en_brightness_export),         // disp_en_brightness.export
		.system_status_export      (controller_inst_system_status_bfm_conduit_export),  //      system_status.export
		.command_en_export         (controller_inst_command_en_export),                 //         command_en.export
		.warning_en_export         (controller_inst_warning_en_export),                 //         warning_en.export
		.boost_export              (controller_inst_boost_export),                      //              boost.export
		.afr_export                (controller_inst_afr_export),                        //                afr.export
		.oil_temp_export           (controller_inst_oil_temp_export),                   //           oil_temp.export
		.coolant_temp_export       (controller_inst_coolant_temp_export),               //       coolant_temp.export
		.intake_temp_export        (controller_inst_intake_temp_export),                //        intake_temp.export
		.ign_en_export             (controller_inst_ign_en_export)                      //             ign_en.export
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) controller_inst_clk_bfm (
		.clk (controller_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_conduit_bfm controller_inst_command_tx_bfm (
		.sig_export (controller_inst_command_tx_export)  // conduit.export
	);

	altera_conduit_bfm_0002 controller_inst_command_rx_bfm (
		.sig_export (controller_inst_command_rx_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0002 controller_inst_command_status_bfm (
		.sig_export (controller_inst_command_status_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0003 controller_inst_disp_en_brightness_bfm (
		.sig_export (controller_inst_disp_en_brightness_export)  // conduit.export
	);

	altera_conduit_bfm_0004 controller_inst_system_status_bfm (
		.sig_export (controller_inst_system_status_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0005 controller_inst_command_en_bfm (
		.sig_export (controller_inst_command_en_export)  // conduit.export
	);

	altera_conduit_bfm_0006 controller_inst_warning_en_bfm (
		.sig_export (controller_inst_warning_en_export)  // conduit.export
	);

	altera_conduit_bfm_0007 controller_inst_boost_bfm (
		.sig_export (controller_inst_boost_export)  // conduit.export
	);

	altera_conduit_bfm_0007 controller_inst_afr_bfm (
		.sig_export (controller_inst_afr_export)  // conduit.export
	);

	altera_conduit_bfm_0007 controller_inst_oil_temp_bfm (
		.sig_export (controller_inst_oil_temp_export)  // conduit.export
	);

	altera_conduit_bfm_0007 controller_inst_coolant_temp_bfm (
		.sig_export (controller_inst_coolant_temp_export)  // conduit.export
	);

	altera_conduit_bfm_0007 controller_inst_intake_temp_bfm (
		.sig_export (controller_inst_intake_temp_export)  // conduit.export
	);

	altera_conduit_bfm_0008 controller_inst_ign_en_bfm (
		.sig_export (controller_inst_ign_en_export)  // conduit.export
	);

endmodule
