// controller_tb.v

// Generated using ACDS version 13.1 162 at 2018.07.10.21:09:13

`timescale 1 ps / 1 ps
module controller_tb (
	);

	wire         controller_inst_clk_bfm_clk_clk;                   // controller_inst_clk_bfm:clk -> controller_inst:clk_clk
	wire   [7:0] controller_inst_command_tx_export;                 // controller_inst:command_tx_export -> controller_inst_command_tx_bfm:sig_export
	wire   [0:0] controller_inst_ign_bfm_conduit_export;            // controller_inst_ign_bfm:sig_export -> controller_inst:ign_export
	wire   [7:0] controller_inst_command_rx_bfm_conduit_export;     // controller_inst_command_rx_bfm:sig_export -> controller_inst:command_rx_export
	wire   [7:0] controller_inst_command_status_bfm_conduit_export; // controller_inst_command_status_bfm:sig_export -> controller_inst:command_status_export
	wire         controller_inst_disp_en_export;                    // controller_inst:disp_en_export -> controller_inst_disp_en_bfm:sig_export
	wire   [7:0] controller_inst_disp_brightness_export;            // controller_inst:disp_brightness_export -> controller_inst_disp_brightness_bfm:sig_export
	wire   [0:0] controller_inst_daylight_bfm_conduit_export;       // controller_inst_daylight_bfm:sig_export -> controller_inst:daylight_export
	wire         controller_inst_conn_export;                       // controller_inst:conn_export -> controller_inst_conn_bfm:sig_export
	wire         controller_inst_err_export;                        // controller_inst:err_export -> controller_inst_err_bfm:sig_export
	wire         controller_inst_command_tx_en_export;              // controller_inst:command_tx_en_export -> controller_inst_command_tx_en_bfm:sig_export
	wire         controller_inst_command_rx_en_export;              // controller_inst:command_rx_en_export -> controller_inst_command_rx_en_bfm:sig_export
	wire         controller_inst_boost_wrn_export;                  // controller_inst:boost_wrn_export -> controller_inst_boost_wrn_bfm:sig_export
	wire         controller_inst_afr_wrn_export;                    // controller_inst:afr_wrn_export -> controller_inst_afr_wrn_bfm:sig_export
	wire         controller_inst_wrn_export;                        // controller_inst:wrn_export -> controller_inst_wrn_bfm:sig_export
	wire  [11:0] controller_inst_boost_export;                      // controller_inst:boost_export -> controller_inst_boost_bfm:sig_export
	wire  [11:0] controller_inst_afr_export;                        // controller_inst:afr_export -> controller_inst_afr_bfm:sig_export
	wire  [11:0] controller_inst_oil_temp_export;                   // controller_inst:oil_temp_export -> controller_inst_oil_temp_bfm:sig_export
	wire  [11:0] controller_inst_coolant_temp_export;               // controller_inst:coolant_temp_export -> controller_inst_coolant_temp_bfm:sig_export
	wire  [11:0] controller_inst_intake_temp_export;                // controller_inst:intake_temp_export -> controller_inst_intake_temp_bfm:sig_export

	controller controller_inst (
		.clk_clk                (controller_inst_clk_bfm_clk_clk),                   //             clk.clk
		.command_tx_export      (controller_inst_command_tx_export),                 //      command_tx.export
		.ign_export             (controller_inst_ign_bfm_conduit_export),            //             ign.export
		.command_rx_export      (controller_inst_command_rx_bfm_conduit_export),     //      command_rx.export
		.command_status_export  (controller_inst_command_status_bfm_conduit_export), //  command_status.export
		.disp_en_export         (controller_inst_disp_en_export),                    //         disp_en.export
		.disp_brightness_export (controller_inst_disp_brightness_export),            // disp_brightness.export
		.daylight_export        (controller_inst_daylight_bfm_conduit_export),       //        daylight.export
		.conn_export            (controller_inst_conn_export),                       //            conn.export
		.err_export             (controller_inst_err_export),                        //             err.export
		.command_tx_en_export   (controller_inst_command_tx_en_export),              //   command_tx_en.export
		.command_rx_en_export   (controller_inst_command_rx_en_export),              //   command_rx_en.export
		.boost_wrn_export       (controller_inst_boost_wrn_export),                  //       boost_wrn.export
		.afr_wrn_export         (controller_inst_afr_wrn_export),                    //         afr_wrn.export
		.wrn_export             (controller_inst_wrn_export),                        //             wrn.export
		.boost_export           (controller_inst_boost_export),                      //           boost.export
		.afr_export             (controller_inst_afr_export),                        //             afr.export
		.oil_temp_export        (controller_inst_oil_temp_export),                   //        oil_temp.export
		.coolant_temp_export    (controller_inst_coolant_temp_export),               //    coolant_temp.export
		.intake_temp_export     (controller_inst_intake_temp_export)                 //     intake_temp.export
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) controller_inst_clk_bfm (
		.clk (controller_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_conduit_bfm controller_inst_command_tx_bfm (
		.sig_export (controller_inst_command_tx_export)  // conduit.export
	);

	altera_conduit_bfm_0002 controller_inst_ign_bfm (
		.sig_export (controller_inst_ign_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0003 controller_inst_command_rx_bfm (
		.sig_export (controller_inst_command_rx_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0003 controller_inst_command_status_bfm (
		.sig_export (controller_inst_command_status_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0004 controller_inst_disp_en_bfm (
		.sig_export (controller_inst_disp_en_export)  // conduit.export
	);

	altera_conduit_bfm controller_inst_disp_brightness_bfm (
		.sig_export (controller_inst_disp_brightness_export)  // conduit.export
	);

	altera_conduit_bfm_0002 controller_inst_daylight_bfm (
		.sig_export (controller_inst_daylight_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0004 controller_inst_conn_bfm (
		.sig_export (controller_inst_conn_export)  // conduit.export
	);

	altera_conduit_bfm_0004 controller_inst_err_bfm (
		.sig_export (controller_inst_err_export)  // conduit.export
	);

	altera_conduit_bfm_0004 controller_inst_command_tx_en_bfm (
		.sig_export (controller_inst_command_tx_en_export)  // conduit.export
	);

	altera_conduit_bfm_0004 controller_inst_command_rx_en_bfm (
		.sig_export (controller_inst_command_rx_en_export)  // conduit.export
	);

	altera_conduit_bfm_0004 controller_inst_boost_wrn_bfm (
		.sig_export (controller_inst_boost_wrn_export)  // conduit.export
	);

	altera_conduit_bfm_0004 controller_inst_afr_wrn_bfm (
		.sig_export (controller_inst_afr_wrn_export)  // conduit.export
	);

	altera_conduit_bfm_0004 controller_inst_wrn_bfm (
		.sig_export (controller_inst_wrn_export)  // conduit.export
	);

	altera_conduit_bfm_0005 controller_inst_boost_bfm (
		.sig_export (controller_inst_boost_export)  // conduit.export
	);

	altera_conduit_bfm_0005 controller_inst_afr_bfm (
		.sig_export (controller_inst_afr_export)  // conduit.export
	);

	altera_conduit_bfm_0005 controller_inst_oil_temp_bfm (
		.sig_export (controller_inst_oil_temp_export)  // conduit.export
	);

	altera_conduit_bfm_0005 controller_inst_coolant_temp_bfm (
		.sig_export (controller_inst_coolant_temp_export)  // conduit.export
	);

	altera_conduit_bfm_0005 controller_inst_intake_temp_bfm (
		.sig_export (controller_inst_intake_temp_export)  // conduit.export
	);

endmodule
