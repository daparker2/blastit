// controller.v

// Generated using ACDS version 13.1 162 at 2018.07.10.21:07:17

`timescale 1 ps / 1 ps
module controller (
		input  wire        clk_clk,                //             clk.clk
		output wire [7:0]  command_tx_export,      //      command_tx.export
		input  wire        ign_export,             //             ign.export
		input  wire [7:0]  command_rx_export,      //      command_rx.export
		input  wire [7:0]  command_status_export,  //  command_status.export
		output wire        disp_en_export,         //         disp_en.export
		output wire [7:0]  disp_brightness_export, // disp_brightness.export
		input  wire        daylight_export,        //        daylight.export
		output wire        conn_export,            //            conn.export
		output wire        err_export,             //             err.export
		output wire        command_tx_en_export,   //   command_tx_en.export
		output wire        command_rx_en_export,   //   command_rx_en.export
		output wire        boost_wrn_export,       //       boost_wrn.export
		output wire        afr_wrn_export,         //         afr_wrn.export
		output wire        wrn_export,             //             wrn.export
		output wire [11:0] boost_export,           //           boost.export
		output wire [11:0] afr_export,             //             afr.export
		output wire [11:0] oil_temp_export,        //        oil_temp.export
		output wire [11:0] coolant_temp_export,    //    coolant_temp.export
		output wire [11:0] intake_temp_export      //     intake_temp.export
	);

	wire         nios2_qsys_0_jtag_debug_module_reset_reset;                   // nios2_qsys_0:jtag_debug_module_resetrequest -> [rst_controller:reset_in0, rst_controller:reset_in1]
	wire  [31:0] mm_interconnect_0_command_rx_en_s1_writedata;                 // mm_interconnect_0:command_rx_en_s1_writedata -> command_rx_en:writedata
	wire   [1:0] mm_interconnect_0_command_rx_en_s1_address;                   // mm_interconnect_0:command_rx_en_s1_address -> command_rx_en:address
	wire         mm_interconnect_0_command_rx_en_s1_chipselect;                // mm_interconnect_0:command_rx_en_s1_chipselect -> command_rx_en:chipselect
	wire         mm_interconnect_0_command_rx_en_s1_write;                     // mm_interconnect_0:command_rx_en_s1_write -> command_rx_en:write_n
	wire  [31:0] mm_interconnect_0_command_rx_en_s1_readdata;                  // command_rx_en:readdata -> mm_interconnect_0:command_rx_en_s1_readdata
	wire  [31:0] mm_interconnect_0_boost_s1_writedata;                         // mm_interconnect_0:boost_s1_writedata -> boost:writedata
	wire   [1:0] mm_interconnect_0_boost_s1_address;                           // mm_interconnect_0:boost_s1_address -> boost:address
	wire         mm_interconnect_0_boost_s1_chipselect;                        // mm_interconnect_0:boost_s1_chipselect -> boost:chipselect
	wire         mm_interconnect_0_boost_s1_write;                             // mm_interconnect_0:boost_s1_write -> boost:write_n
	wire  [31:0] mm_interconnect_0_boost_s1_readdata;                          // boost:readdata -> mm_interconnect_0:boost_s1_readdata
	wire         nios2_qsys_0_instruction_master_waitrequest;                  // mm_interconnect_0:nios2_qsys_0_instruction_master_waitrequest -> nios2_qsys_0:i_waitrequest
	wire  [13:0] nios2_qsys_0_instruction_master_address;                      // nios2_qsys_0:i_address -> mm_interconnect_0:nios2_qsys_0_instruction_master_address
	wire         nios2_qsys_0_instruction_master_read;                         // nios2_qsys_0:i_read -> mm_interconnect_0:nios2_qsys_0_instruction_master_read
	wire  [31:0] nios2_qsys_0_instruction_master_readdata;                     // mm_interconnect_0:nios2_qsys_0_instruction_master_readdata -> nios2_qsys_0:i_readdata
	wire         nios2_qsys_0_instruction_master_readdatavalid;                // mm_interconnect_0:nios2_qsys_0_instruction_master_readdatavalid -> nios2_qsys_0:i_readdatavalid
	wire   [0:0] mm_interconnect_0_sysid_c001_control_slave_address;           // mm_interconnect_0:sysid_c001_control_slave_address -> sysid_c001:address
	wire  [31:0] mm_interconnect_0_sysid_c001_control_slave_readdata;          // sysid_c001:readdata -> mm_interconnect_0:sysid_c001_control_slave_readdata
	wire  [31:0] mm_interconnect_0_disp_en_s1_writedata;                       // mm_interconnect_0:disp_en_s1_writedata -> disp_en:writedata
	wire   [1:0] mm_interconnect_0_disp_en_s1_address;                         // mm_interconnect_0:disp_en_s1_address -> disp_en:address
	wire         mm_interconnect_0_disp_en_s1_chipselect;                      // mm_interconnect_0:disp_en_s1_chipselect -> disp_en:chipselect
	wire         mm_interconnect_0_disp_en_s1_write;                           // mm_interconnect_0:disp_en_s1_write -> disp_en:write_n
	wire  [31:0] mm_interconnect_0_disp_en_s1_readdata;                        // disp_en:readdata -> mm_interconnect_0:disp_en_s1_readdata
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest; // nios2_qsys_0:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata;   // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_writedata -> nios2_qsys_0:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address;     // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_address -> nios2_qsys_0:jtag_debug_module_address
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write;       // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_write -> nios2_qsys_0:jtag_debug_module_write
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read;        // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_read -> nios2_qsys_0:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata;    // nios2_qsys_0:jtag_debug_module_readdata -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess; // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_debugaccess -> nios2_qsys_0:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable;  // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_byteenable -> nios2_qsys_0:jtag_debug_module_byteenable
	wire  [31:0] mm_interconnect_0_command_tx_en_s1_writedata;                 // mm_interconnect_0:command_tx_en_s1_writedata -> command_tx_en:writedata
	wire   [1:0] mm_interconnect_0_command_tx_en_s1_address;                   // mm_interconnect_0:command_tx_en_s1_address -> command_tx_en:address
	wire         mm_interconnect_0_command_tx_en_s1_chipselect;                // mm_interconnect_0:command_tx_en_s1_chipselect -> command_tx_en:chipselect
	wire         mm_interconnect_0_command_tx_en_s1_write;                     // mm_interconnect_0:command_tx_en_s1_write -> command_tx_en:write_n
	wire  [31:0] mm_interconnect_0_command_tx_en_s1_readdata;                  // command_tx_en:readdata -> mm_interconnect_0:command_tx_en_s1_readdata
	wire  [31:0] mm_interconnect_0_iram_s1_writedata;                          // mm_interconnect_0:iram_s1_writedata -> iram:writedata
	wire   [8:0] mm_interconnect_0_iram_s1_address;                            // mm_interconnect_0:iram_s1_address -> iram:address
	wire         mm_interconnect_0_iram_s1_chipselect;                         // mm_interconnect_0:iram_s1_chipselect -> iram:chipselect
	wire         mm_interconnect_0_iram_s1_clken;                              // mm_interconnect_0:iram_s1_clken -> iram:clken
	wire         mm_interconnect_0_iram_s1_write;                              // mm_interconnect_0:iram_s1_write -> iram:write
	wire  [31:0] mm_interconnect_0_iram_s1_readdata;                           // iram:readdata -> mm_interconnect_0:iram_s1_readdata
	wire         mm_interconnect_0_iram_s1_debugaccess;                        // mm_interconnect_0:iram_s1_debugaccess -> iram:debugaccess
	wire   [3:0] mm_interconnect_0_iram_s1_byteenable;                         // mm_interconnect_0:iram_s1_byteenable -> iram:byteenable
	wire   [1:0] mm_interconnect_0_daylight_s1_address;                        // mm_interconnect_0:daylight_s1_address -> daylight:address
	wire  [31:0] mm_interconnect_0_daylight_s1_readdata;                       // daylight:readdata -> mm_interconnect_0:daylight_s1_readdata
	wire  [31:0] mm_interconnect_0_command_tx_s1_writedata;                    // mm_interconnect_0:command_tx_s1_writedata -> command_tx:writedata
	wire   [1:0] mm_interconnect_0_command_tx_s1_address;                      // mm_interconnect_0:command_tx_s1_address -> command_tx:address
	wire         mm_interconnect_0_command_tx_s1_chipselect;                   // mm_interconnect_0:command_tx_s1_chipselect -> command_tx:chipselect
	wire         mm_interconnect_0_command_tx_s1_write;                        // mm_interconnect_0:command_tx_s1_write -> command_tx:write_n
	wire  [31:0] mm_interconnect_0_command_tx_s1_readdata;                     // command_tx:readdata -> mm_interconnect_0:command_tx_s1_readdata
	wire   [1:0] mm_interconnect_0_ign_s1_address;                             // mm_interconnect_0:ign_s1_address -> ign:address
	wire  [31:0] mm_interconnect_0_ign_s1_readdata;                            // ign:readdata -> mm_interconnect_0:ign_s1_readdata
	wire  [31:0] mm_interconnect_0_afr_wrn_s1_writedata;                       // mm_interconnect_0:afr_wrn_s1_writedata -> afr_wrn:writedata
	wire   [1:0] mm_interconnect_0_afr_wrn_s1_address;                         // mm_interconnect_0:afr_wrn_s1_address -> afr_wrn:address
	wire         mm_interconnect_0_afr_wrn_s1_chipselect;                      // mm_interconnect_0:afr_wrn_s1_chipselect -> afr_wrn:chipselect
	wire         mm_interconnect_0_afr_wrn_s1_write;                           // mm_interconnect_0:afr_wrn_s1_write -> afr_wrn:write_n
	wire  [31:0] mm_interconnect_0_afr_wrn_s1_readdata;                        // afr_wrn:readdata -> mm_interconnect_0:afr_wrn_s1_readdata
	wire   [1:0] mm_interconnect_0_command_status_s1_address;                  // mm_interconnect_0:command_status_s1_address -> command_status:address
	wire  [31:0] mm_interconnect_0_command_status_s1_readdata;                 // command_status:readdata -> mm_interconnect_0:command_status_s1_readdata
	wire  [31:0] mm_interconnect_0_boost_wrn_s1_writedata;                     // mm_interconnect_0:boost_wrn_s1_writedata -> boost_wrn:writedata
	wire   [1:0] mm_interconnect_0_boost_wrn_s1_address;                       // mm_interconnect_0:boost_wrn_s1_address -> boost_wrn:address
	wire         mm_interconnect_0_boost_wrn_s1_chipselect;                    // mm_interconnect_0:boost_wrn_s1_chipselect -> boost_wrn:chipselect
	wire         mm_interconnect_0_boost_wrn_s1_write;                         // mm_interconnect_0:boost_wrn_s1_write -> boost_wrn:write_n
	wire  [31:0] mm_interconnect_0_boost_wrn_s1_readdata;                      // boost_wrn:readdata -> mm_interconnect_0:boost_wrn_s1_readdata
	wire  [31:0] mm_interconnect_0_intake_temp_s1_writedata;                   // mm_interconnect_0:intake_temp_s1_writedata -> intake_temp:writedata
	wire   [1:0] mm_interconnect_0_intake_temp_s1_address;                     // mm_interconnect_0:intake_temp_s1_address -> intake_temp:address
	wire         mm_interconnect_0_intake_temp_s1_chipselect;                  // mm_interconnect_0:intake_temp_s1_chipselect -> intake_temp:chipselect
	wire         mm_interconnect_0_intake_temp_s1_write;                       // mm_interconnect_0:intake_temp_s1_write -> intake_temp:write_n
	wire  [31:0] mm_interconnect_0_intake_temp_s1_readdata;                    // intake_temp:readdata -> mm_interconnect_0:intake_temp_s1_readdata
	wire  [31:0] mm_interconnect_0_err_s1_writedata;                           // mm_interconnect_0:err_s1_writedata -> err:writedata
	wire   [1:0] mm_interconnect_0_err_s1_address;                             // mm_interconnect_0:err_s1_address -> err:address
	wire         mm_interconnect_0_err_s1_chipselect;                          // mm_interconnect_0:err_s1_chipselect -> err:chipselect
	wire         mm_interconnect_0_err_s1_write;                               // mm_interconnect_0:err_s1_write -> err:write_n
	wire  [31:0] mm_interconnect_0_err_s1_readdata;                            // err:readdata -> mm_interconnect_0:err_s1_readdata
	wire   [1:0] mm_interconnect_0_command_rx_s1_address;                      // mm_interconnect_0:command_rx_s1_address -> command_rx:address
	wire  [31:0] mm_interconnect_0_command_rx_s1_readdata;                     // command_rx:readdata -> mm_interconnect_0:command_rx_s1_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;  // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;    // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;      // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;         // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;     // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire  [31:0] mm_interconnect_0_wrn_s1_writedata;                           // mm_interconnect_0:wrn_s1_writedata -> wrn:writedata
	wire   [1:0] mm_interconnect_0_wrn_s1_address;                             // mm_interconnect_0:wrn_s1_address -> wrn:address
	wire         mm_interconnect_0_wrn_s1_chipselect;                          // mm_interconnect_0:wrn_s1_chipselect -> wrn:chipselect
	wire         mm_interconnect_0_wrn_s1_write;                               // mm_interconnect_0:wrn_s1_write -> wrn:write_n
	wire  [31:0] mm_interconnect_0_wrn_s1_readdata;                            // wrn:readdata -> mm_interconnect_0:wrn_s1_readdata
	wire  [31:0] mm_interconnect_0_disp_brightness_s1_writedata;               // mm_interconnect_0:disp_brightness_s1_writedata -> disp_brightness:writedata
	wire   [1:0] mm_interconnect_0_disp_brightness_s1_address;                 // mm_interconnect_0:disp_brightness_s1_address -> disp_brightness:address
	wire         mm_interconnect_0_disp_brightness_s1_chipselect;              // mm_interconnect_0:disp_brightness_s1_chipselect -> disp_brightness:chipselect
	wire         mm_interconnect_0_disp_brightness_s1_write;                   // mm_interconnect_0:disp_brightness_s1_write -> disp_brightness:write_n
	wire  [31:0] mm_interconnect_0_disp_brightness_s1_readdata;                // disp_brightness:readdata -> mm_interconnect_0:disp_brightness_s1_readdata
	wire  [31:0] mm_interconnect_0_conn_s1_writedata;                          // mm_interconnect_0:conn_s1_writedata -> conn:writedata
	wire   [1:0] mm_interconnect_0_conn_s1_address;                            // mm_interconnect_0:conn_s1_address -> conn:address
	wire         mm_interconnect_0_conn_s1_chipselect;                         // mm_interconnect_0:conn_s1_chipselect -> conn:chipselect
	wire         mm_interconnect_0_conn_s1_write;                              // mm_interconnect_0:conn_s1_write -> conn:write_n
	wire  [31:0] mm_interconnect_0_conn_s1_readdata;                           // conn:readdata -> mm_interconnect_0:conn_s1_readdata
	wire  [31:0] mm_interconnect_0_dram_s1_writedata;                          // mm_interconnect_0:dram_s1_writedata -> dram:writedata
	wire   [8:0] mm_interconnect_0_dram_s1_address;                            // mm_interconnect_0:dram_s1_address -> dram:address
	wire         mm_interconnect_0_dram_s1_chipselect;                         // mm_interconnect_0:dram_s1_chipselect -> dram:chipselect
	wire         mm_interconnect_0_dram_s1_clken;                              // mm_interconnect_0:dram_s1_clken -> dram:clken
	wire         mm_interconnect_0_dram_s1_write;                              // mm_interconnect_0:dram_s1_write -> dram:write
	wire  [31:0] mm_interconnect_0_dram_s1_readdata;                           // dram:readdata -> mm_interconnect_0:dram_s1_readdata
	wire   [3:0] mm_interconnect_0_dram_s1_byteenable;                         // mm_interconnect_0:dram_s1_byteenable -> dram:byteenable
	wire  [31:0] mm_interconnect_0_afr_s1_writedata;                           // mm_interconnect_0:afr_s1_writedata -> afr:writedata
	wire   [1:0] mm_interconnect_0_afr_s1_address;                             // mm_interconnect_0:afr_s1_address -> afr:address
	wire         mm_interconnect_0_afr_s1_chipselect;                          // mm_interconnect_0:afr_s1_chipselect -> afr:chipselect
	wire         mm_interconnect_0_afr_s1_write;                               // mm_interconnect_0:afr_s1_write -> afr:write_n
	wire  [31:0] mm_interconnect_0_afr_s1_readdata;                            // afr:readdata -> mm_interconnect_0:afr_s1_readdata
	wire  [31:0] mm_interconnect_0_coolant_temp_s1_writedata;                  // mm_interconnect_0:coolant_temp_s1_writedata -> coolant_temp:writedata
	wire   [1:0] mm_interconnect_0_coolant_temp_s1_address;                    // mm_interconnect_0:coolant_temp_s1_address -> coolant_temp:address
	wire         mm_interconnect_0_coolant_temp_s1_chipselect;                 // mm_interconnect_0:coolant_temp_s1_chipselect -> coolant_temp:chipselect
	wire         mm_interconnect_0_coolant_temp_s1_write;                      // mm_interconnect_0:coolant_temp_s1_write -> coolant_temp:write_n
	wire  [31:0] mm_interconnect_0_coolant_temp_s1_readdata;                   // coolant_temp:readdata -> mm_interconnect_0:coolant_temp_s1_readdata
	wire  [31:0] mm_interconnect_0_oil_temp_s1_writedata;                      // mm_interconnect_0:oil_temp_s1_writedata -> oil_temp:writedata
	wire   [1:0] mm_interconnect_0_oil_temp_s1_address;                        // mm_interconnect_0:oil_temp_s1_address -> oil_temp:address
	wire         mm_interconnect_0_oil_temp_s1_chipselect;                     // mm_interconnect_0:oil_temp_s1_chipselect -> oil_temp:chipselect
	wire         mm_interconnect_0_oil_temp_s1_write;                          // mm_interconnect_0:oil_temp_s1_write -> oil_temp:write_n
	wire  [31:0] mm_interconnect_0_oil_temp_s1_readdata;                       // oil_temp:readdata -> mm_interconnect_0:oil_temp_s1_readdata
	wire         nios2_qsys_0_data_master_waitrequest;                         // mm_interconnect_0:nios2_qsys_0_data_master_waitrequest -> nios2_qsys_0:d_waitrequest
	wire  [31:0] nios2_qsys_0_data_master_writedata;                           // nios2_qsys_0:d_writedata -> mm_interconnect_0:nios2_qsys_0_data_master_writedata
	wire  [13:0] nios2_qsys_0_data_master_address;                             // nios2_qsys_0:d_address -> mm_interconnect_0:nios2_qsys_0_data_master_address
	wire         nios2_qsys_0_data_master_write;                               // nios2_qsys_0:d_write -> mm_interconnect_0:nios2_qsys_0_data_master_write
	wire         nios2_qsys_0_data_master_read;                                // nios2_qsys_0:d_read -> mm_interconnect_0:nios2_qsys_0_data_master_read
	wire  [31:0] nios2_qsys_0_data_master_readdata;                            // mm_interconnect_0:nios2_qsys_0_data_master_readdata -> nios2_qsys_0:d_readdata
	wire         nios2_qsys_0_data_master_debugaccess;                         // nios2_qsys_0:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_0_data_master_debugaccess
	wire         nios2_qsys_0_data_master_readdatavalid;                       // mm_interconnect_0:nios2_qsys_0_data_master_readdatavalid -> nios2_qsys_0:d_readdatavalid
	wire   [3:0] nios2_qsys_0_data_master_byteenable;                          // nios2_qsys_0:d_byteenable -> mm_interconnect_0:nios2_qsys_0_data_master_byteenable
	wire         irq_mapper_receiver0_irq;                                     // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_qsys_0_d_irq_irq;                                       // irq_mapper:sender_irq -> nios2_qsys_0:d_irq
	wire         rst_controller_reset_out_reset;                               // rst_controller:reset_out -> [afr:reset_n, afr_wrn:reset_n, boost:reset_n, boost_wrn:reset_n, command_rx:reset_n, command_rx_en:reset_n, command_status:reset_n, command_tx:reset_n, command_tx_en:reset_n, conn:reset_n, coolant_temp:reset_n, daylight:reset_n, disp_brightness:reset_n, disp_en:reset_n, dram:reset, err:reset_n, ign:reset_n, intake_temp:reset_n, iram:reset, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:nios2_qsys_0_reset_n_reset_bridge_in_reset_reset, nios2_qsys_0:reset_n, oil_temp:reset_n, rst_translator:in_reset, sysid_c001:reset_n, wrn:reset_n]
	wire         rst_controller_reset_out_reset_req;                           // rst_controller:reset_req -> [dram:reset_req, iram:reset_req, nios2_qsys_0:reset_req, rst_translator:reset_req_in]

	controller_nios2_qsys_0 nios2_qsys_0 (
		.clk                                   (clk_clk),                                                      //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                              //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                           //                          .reset_req
		.d_address                             (nios2_qsys_0_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_qsys_0_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_qsys_0_data_master_read),                                //                          .read
		.d_readdata                            (nios2_qsys_0_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_qsys_0_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_qsys_0_data_master_write),                               //                          .write
		.d_writedata                           (nios2_qsys_0_data_master_writedata),                           //                          .writedata
		.d_readdatavalid                       (nios2_qsys_0_data_master_readdatavalid),                       //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_0_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_qsys_0_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_qsys_0_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_qsys_0_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_qsys_0_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (nios2_qsys_0_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (nios2_qsys_0_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_qsys_0_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                              // custom_instruction_master.readra
	);

	controller_dram dram (
		.clk        (clk_clk),                              //   clk1.clk
		.address    (mm_interconnect_0_dram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_dram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_dram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_dram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_dram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_dram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_dram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),       // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)    //       .reset_req
	);

	controller_sysid_c001 sysid_c001 (
		.clock    (clk_clk),                                             //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                     //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_c001_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_c001_control_slave_address)   //              .address
	);

	controller_iram iram (
		.clk         (clk_clk),                               //   clk1.clk
		.address     (mm_interconnect_0_iram_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_iram_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_iram_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_iram_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_iram_s1_write),       //       .write
		.readdata    (mm_interconnect_0_iram_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_iram_s1_writedata),   //       .writedata
		.byteenable  (mm_interconnect_0_iram_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),        // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req)     //       .reset_req
	);

	controller_ign ign (
		.clk      (clk_clk),                           //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),   //               reset.reset_n
		.address  (mm_interconnect_0_ign_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_ign_s1_readdata), //                    .readdata
		.in_port  (ign_export)                         // external_connection.export
	);

	controller_command_tx command_tx (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_command_tx_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_command_tx_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_command_tx_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_command_tx_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_command_tx_s1_readdata),   //                    .readdata
		.out_port   (command_tx_export)                           // external_connection.export
	);

	controller_command_rx command_rx (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_command_rx_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_command_rx_s1_readdata), //                    .readdata
		.in_port  (command_rx_export)                         // external_connection.export
	);

	controller_command_rx command_status (
		.clk      (clk_clk),                                      //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address  (mm_interconnect_0_command_status_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_command_status_s1_readdata), //                    .readdata
		.in_port  (command_status_export)                         // external_connection.export
	);

	controller_disp_en disp_en (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_disp_en_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_disp_en_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_disp_en_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_disp_en_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_disp_en_s1_readdata),   //                    .readdata
		.out_port   (disp_en_export)                           // external_connection.export
	);

	controller_command_tx disp_brightness (
		.clk        (clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_disp_brightness_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_disp_brightness_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_disp_brightness_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_disp_brightness_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_disp_brightness_s1_readdata),   //                    .readdata
		.out_port   (disp_brightness_export)                           // external_connection.export
	);

	controller_ign daylight (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_daylight_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_daylight_s1_readdata), //                    .readdata
		.in_port  (daylight_export)                         // external_connection.export
	);

	controller_disp_en conn (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_conn_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_conn_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_conn_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_conn_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_conn_s1_readdata),   //                    .readdata
		.out_port   (conn_export)                           // external_connection.export
	);

	controller_disp_en err (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_err_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_err_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_err_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_err_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_err_s1_readdata),   //                    .readdata
		.out_port   (err_export)                           // external_connection.export
	);

	controller_disp_en command_tx_en (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_command_tx_en_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_command_tx_en_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_command_tx_en_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_command_tx_en_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_command_tx_en_s1_readdata),   //                    .readdata
		.out_port   (command_tx_en_export)                           // external_connection.export
	);

	controller_disp_en command_rx_en (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_command_rx_en_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_command_rx_en_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_command_rx_en_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_command_rx_en_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_command_rx_en_s1_readdata),   //                    .readdata
		.out_port   (command_rx_en_export)                           // external_connection.export
	);

	controller_disp_en boost_wrn (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_boost_wrn_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_boost_wrn_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_boost_wrn_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_boost_wrn_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_boost_wrn_s1_readdata),   //                    .readdata
		.out_port   (boost_wrn_export)                           // external_connection.export
	);

	controller_disp_en afr_wrn (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_afr_wrn_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_afr_wrn_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_afr_wrn_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_afr_wrn_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_afr_wrn_s1_readdata),   //                    .readdata
		.out_port   (afr_wrn_export)                           // external_connection.export
	);

	controller_disp_en wrn (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_wrn_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_wrn_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_wrn_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_wrn_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_wrn_s1_readdata),   //                    .readdata
		.out_port   (wrn_export)                           // external_connection.export
	);

	controller_boost boost (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_boost_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_boost_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_boost_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_boost_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_boost_s1_readdata),   //                    .readdata
		.out_port   (boost_export)                           // external_connection.export
	);

	controller_boost afr (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_afr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_afr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_afr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_afr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_afr_s1_readdata),   //                    .readdata
		.out_port   (afr_export)                           // external_connection.export
	);

	controller_boost oil_temp (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_oil_temp_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_oil_temp_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_oil_temp_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_oil_temp_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_oil_temp_s1_readdata),   //                    .readdata
		.out_port   (oil_temp_export)                           // external_connection.export
	);

	controller_boost coolant_temp (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_coolant_temp_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_coolant_temp_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_coolant_temp_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_coolant_temp_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_coolant_temp_s1_readdata),   //                    .readdata
		.out_port   (coolant_temp_export)                           // external_connection.export
	);

	controller_boost intake_temp (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_intake_temp_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_intake_temp_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_intake_temp_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_intake_temp_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_intake_temp_s1_readdata),   //                    .readdata
		.out_port   (intake_temp_export)                           // external_connection.export
	);

	controller_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	controller_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                    (clk_clk),                                                      //                                  clk_0_clk.clk
		.nios2_qsys_0_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                               // nios2_qsys_0_reset_n_reset_bridge_in_reset.reset
		.nios2_qsys_0_data_master_address                 (nios2_qsys_0_data_master_address),                             //                   nios2_qsys_0_data_master.address
		.nios2_qsys_0_data_master_waitrequest             (nios2_qsys_0_data_master_waitrequest),                         //                                           .waitrequest
		.nios2_qsys_0_data_master_byteenable              (nios2_qsys_0_data_master_byteenable),                          //                                           .byteenable
		.nios2_qsys_0_data_master_read                    (nios2_qsys_0_data_master_read),                                //                                           .read
		.nios2_qsys_0_data_master_readdata                (nios2_qsys_0_data_master_readdata),                            //                                           .readdata
		.nios2_qsys_0_data_master_readdatavalid           (nios2_qsys_0_data_master_readdatavalid),                       //                                           .readdatavalid
		.nios2_qsys_0_data_master_write                   (nios2_qsys_0_data_master_write),                               //                                           .write
		.nios2_qsys_0_data_master_writedata               (nios2_qsys_0_data_master_writedata),                           //                                           .writedata
		.nios2_qsys_0_data_master_debugaccess             (nios2_qsys_0_data_master_debugaccess),                         //                                           .debugaccess
		.nios2_qsys_0_instruction_master_address          (nios2_qsys_0_instruction_master_address),                      //            nios2_qsys_0_instruction_master.address
		.nios2_qsys_0_instruction_master_waitrequest      (nios2_qsys_0_instruction_master_waitrequest),                  //                                           .waitrequest
		.nios2_qsys_0_instruction_master_read             (nios2_qsys_0_instruction_master_read),                         //                                           .read
		.nios2_qsys_0_instruction_master_readdata         (nios2_qsys_0_instruction_master_readdata),                     //                                           .readdata
		.nios2_qsys_0_instruction_master_readdatavalid    (nios2_qsys_0_instruction_master_readdatavalid),                //                                           .readdatavalid
		.afr_s1_address                                   (mm_interconnect_0_afr_s1_address),                             //                                     afr_s1.address
		.afr_s1_write                                     (mm_interconnect_0_afr_s1_write),                               //                                           .write
		.afr_s1_readdata                                  (mm_interconnect_0_afr_s1_readdata),                            //                                           .readdata
		.afr_s1_writedata                                 (mm_interconnect_0_afr_s1_writedata),                           //                                           .writedata
		.afr_s1_chipselect                                (mm_interconnect_0_afr_s1_chipselect),                          //                                           .chipselect
		.afr_wrn_s1_address                               (mm_interconnect_0_afr_wrn_s1_address),                         //                                 afr_wrn_s1.address
		.afr_wrn_s1_write                                 (mm_interconnect_0_afr_wrn_s1_write),                           //                                           .write
		.afr_wrn_s1_readdata                              (mm_interconnect_0_afr_wrn_s1_readdata),                        //                                           .readdata
		.afr_wrn_s1_writedata                             (mm_interconnect_0_afr_wrn_s1_writedata),                       //                                           .writedata
		.afr_wrn_s1_chipselect                            (mm_interconnect_0_afr_wrn_s1_chipselect),                      //                                           .chipselect
		.boost_s1_address                                 (mm_interconnect_0_boost_s1_address),                           //                                   boost_s1.address
		.boost_s1_write                                   (mm_interconnect_0_boost_s1_write),                             //                                           .write
		.boost_s1_readdata                                (mm_interconnect_0_boost_s1_readdata),                          //                                           .readdata
		.boost_s1_writedata                               (mm_interconnect_0_boost_s1_writedata),                         //                                           .writedata
		.boost_s1_chipselect                              (mm_interconnect_0_boost_s1_chipselect),                        //                                           .chipselect
		.boost_wrn_s1_address                             (mm_interconnect_0_boost_wrn_s1_address),                       //                               boost_wrn_s1.address
		.boost_wrn_s1_write                               (mm_interconnect_0_boost_wrn_s1_write),                         //                                           .write
		.boost_wrn_s1_readdata                            (mm_interconnect_0_boost_wrn_s1_readdata),                      //                                           .readdata
		.boost_wrn_s1_writedata                           (mm_interconnect_0_boost_wrn_s1_writedata),                     //                                           .writedata
		.boost_wrn_s1_chipselect                          (mm_interconnect_0_boost_wrn_s1_chipselect),                    //                                           .chipselect
		.command_rx_s1_address                            (mm_interconnect_0_command_rx_s1_address),                      //                              command_rx_s1.address
		.command_rx_s1_readdata                           (mm_interconnect_0_command_rx_s1_readdata),                     //                                           .readdata
		.command_rx_en_s1_address                         (mm_interconnect_0_command_rx_en_s1_address),                   //                           command_rx_en_s1.address
		.command_rx_en_s1_write                           (mm_interconnect_0_command_rx_en_s1_write),                     //                                           .write
		.command_rx_en_s1_readdata                        (mm_interconnect_0_command_rx_en_s1_readdata),                  //                                           .readdata
		.command_rx_en_s1_writedata                       (mm_interconnect_0_command_rx_en_s1_writedata),                 //                                           .writedata
		.command_rx_en_s1_chipselect                      (mm_interconnect_0_command_rx_en_s1_chipselect),                //                                           .chipselect
		.command_status_s1_address                        (mm_interconnect_0_command_status_s1_address),                  //                          command_status_s1.address
		.command_status_s1_readdata                       (mm_interconnect_0_command_status_s1_readdata),                 //                                           .readdata
		.command_tx_s1_address                            (mm_interconnect_0_command_tx_s1_address),                      //                              command_tx_s1.address
		.command_tx_s1_write                              (mm_interconnect_0_command_tx_s1_write),                        //                                           .write
		.command_tx_s1_readdata                           (mm_interconnect_0_command_tx_s1_readdata),                     //                                           .readdata
		.command_tx_s1_writedata                          (mm_interconnect_0_command_tx_s1_writedata),                    //                                           .writedata
		.command_tx_s1_chipselect                         (mm_interconnect_0_command_tx_s1_chipselect),                   //                                           .chipselect
		.command_tx_en_s1_address                         (mm_interconnect_0_command_tx_en_s1_address),                   //                           command_tx_en_s1.address
		.command_tx_en_s1_write                           (mm_interconnect_0_command_tx_en_s1_write),                     //                                           .write
		.command_tx_en_s1_readdata                        (mm_interconnect_0_command_tx_en_s1_readdata),                  //                                           .readdata
		.command_tx_en_s1_writedata                       (mm_interconnect_0_command_tx_en_s1_writedata),                 //                                           .writedata
		.command_tx_en_s1_chipselect                      (mm_interconnect_0_command_tx_en_s1_chipselect),                //                                           .chipselect
		.conn_s1_address                                  (mm_interconnect_0_conn_s1_address),                            //                                    conn_s1.address
		.conn_s1_write                                    (mm_interconnect_0_conn_s1_write),                              //                                           .write
		.conn_s1_readdata                                 (mm_interconnect_0_conn_s1_readdata),                           //                                           .readdata
		.conn_s1_writedata                                (mm_interconnect_0_conn_s1_writedata),                          //                                           .writedata
		.conn_s1_chipselect                               (mm_interconnect_0_conn_s1_chipselect),                         //                                           .chipselect
		.coolant_temp_s1_address                          (mm_interconnect_0_coolant_temp_s1_address),                    //                            coolant_temp_s1.address
		.coolant_temp_s1_write                            (mm_interconnect_0_coolant_temp_s1_write),                      //                                           .write
		.coolant_temp_s1_readdata                         (mm_interconnect_0_coolant_temp_s1_readdata),                   //                                           .readdata
		.coolant_temp_s1_writedata                        (mm_interconnect_0_coolant_temp_s1_writedata),                  //                                           .writedata
		.coolant_temp_s1_chipselect                       (mm_interconnect_0_coolant_temp_s1_chipselect),                 //                                           .chipselect
		.daylight_s1_address                              (mm_interconnect_0_daylight_s1_address),                        //                                daylight_s1.address
		.daylight_s1_readdata                             (mm_interconnect_0_daylight_s1_readdata),                       //                                           .readdata
		.disp_brightness_s1_address                       (mm_interconnect_0_disp_brightness_s1_address),                 //                         disp_brightness_s1.address
		.disp_brightness_s1_write                         (mm_interconnect_0_disp_brightness_s1_write),                   //                                           .write
		.disp_brightness_s1_readdata                      (mm_interconnect_0_disp_brightness_s1_readdata),                //                                           .readdata
		.disp_brightness_s1_writedata                     (mm_interconnect_0_disp_brightness_s1_writedata),               //                                           .writedata
		.disp_brightness_s1_chipselect                    (mm_interconnect_0_disp_brightness_s1_chipselect),              //                                           .chipselect
		.disp_en_s1_address                               (mm_interconnect_0_disp_en_s1_address),                         //                                 disp_en_s1.address
		.disp_en_s1_write                                 (mm_interconnect_0_disp_en_s1_write),                           //                                           .write
		.disp_en_s1_readdata                              (mm_interconnect_0_disp_en_s1_readdata),                        //                                           .readdata
		.disp_en_s1_writedata                             (mm_interconnect_0_disp_en_s1_writedata),                       //                                           .writedata
		.disp_en_s1_chipselect                            (mm_interconnect_0_disp_en_s1_chipselect),                      //                                           .chipselect
		.dram_s1_address                                  (mm_interconnect_0_dram_s1_address),                            //                                    dram_s1.address
		.dram_s1_write                                    (mm_interconnect_0_dram_s1_write),                              //                                           .write
		.dram_s1_readdata                                 (mm_interconnect_0_dram_s1_readdata),                           //                                           .readdata
		.dram_s1_writedata                                (mm_interconnect_0_dram_s1_writedata),                          //                                           .writedata
		.dram_s1_byteenable                               (mm_interconnect_0_dram_s1_byteenable),                         //                                           .byteenable
		.dram_s1_chipselect                               (mm_interconnect_0_dram_s1_chipselect),                         //                                           .chipselect
		.dram_s1_clken                                    (mm_interconnect_0_dram_s1_clken),                              //                                           .clken
		.err_s1_address                                   (mm_interconnect_0_err_s1_address),                             //                                     err_s1.address
		.err_s1_write                                     (mm_interconnect_0_err_s1_write),                               //                                           .write
		.err_s1_readdata                                  (mm_interconnect_0_err_s1_readdata),                            //                                           .readdata
		.err_s1_writedata                                 (mm_interconnect_0_err_s1_writedata),                           //                                           .writedata
		.err_s1_chipselect                                (mm_interconnect_0_err_s1_chipselect),                          //                                           .chipselect
		.ign_s1_address                                   (mm_interconnect_0_ign_s1_address),                             //                                     ign_s1.address
		.ign_s1_readdata                                  (mm_interconnect_0_ign_s1_readdata),                            //                                           .readdata
		.intake_temp_s1_address                           (mm_interconnect_0_intake_temp_s1_address),                     //                             intake_temp_s1.address
		.intake_temp_s1_write                             (mm_interconnect_0_intake_temp_s1_write),                       //                                           .write
		.intake_temp_s1_readdata                          (mm_interconnect_0_intake_temp_s1_readdata),                    //                                           .readdata
		.intake_temp_s1_writedata                         (mm_interconnect_0_intake_temp_s1_writedata),                   //                                           .writedata
		.intake_temp_s1_chipselect                        (mm_interconnect_0_intake_temp_s1_chipselect),                  //                                           .chipselect
		.iram_s1_address                                  (mm_interconnect_0_iram_s1_address),                            //                                    iram_s1.address
		.iram_s1_write                                    (mm_interconnect_0_iram_s1_write),                              //                                           .write
		.iram_s1_readdata                                 (mm_interconnect_0_iram_s1_readdata),                           //                                           .readdata
		.iram_s1_writedata                                (mm_interconnect_0_iram_s1_writedata),                          //                                           .writedata
		.iram_s1_byteenable                               (mm_interconnect_0_iram_s1_byteenable),                         //                                           .byteenable
		.iram_s1_chipselect                               (mm_interconnect_0_iram_s1_chipselect),                         //                                           .chipselect
		.iram_s1_clken                                    (mm_interconnect_0_iram_s1_clken),                              //                                           .clken
		.iram_s1_debugaccess                              (mm_interconnect_0_iram_s1_debugaccess),                        //                                           .debugaccess
		.jtag_uart_0_avalon_jtag_slave_address            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),      //              jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write              (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),        //                                           .write
		.jtag_uart_0_avalon_jtag_slave_read               (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),         //                                           .read
		.jtag_uart_0_avalon_jtag_slave_readdata           (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),     //                                           .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),    //                                           .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),  //                                           .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),   //                                           .chipselect
		.nios2_qsys_0_jtag_debug_module_address           (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),     //             nios2_qsys_0_jtag_debug_module.address
		.nios2_qsys_0_jtag_debug_module_write             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),       //                                           .write
		.nios2_qsys_0_jtag_debug_module_read              (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),        //                                           .read
		.nios2_qsys_0_jtag_debug_module_readdata          (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),    //                                           .readdata
		.nios2_qsys_0_jtag_debug_module_writedata         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),   //                                           .writedata
		.nios2_qsys_0_jtag_debug_module_byteenable        (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),  //                                           .byteenable
		.nios2_qsys_0_jtag_debug_module_waitrequest       (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest), //                                           .waitrequest
		.nios2_qsys_0_jtag_debug_module_debugaccess       (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess), //                                           .debugaccess
		.oil_temp_s1_address                              (mm_interconnect_0_oil_temp_s1_address),                        //                                oil_temp_s1.address
		.oil_temp_s1_write                                (mm_interconnect_0_oil_temp_s1_write),                          //                                           .write
		.oil_temp_s1_readdata                             (mm_interconnect_0_oil_temp_s1_readdata),                       //                                           .readdata
		.oil_temp_s1_writedata                            (mm_interconnect_0_oil_temp_s1_writedata),                      //                                           .writedata
		.oil_temp_s1_chipselect                           (mm_interconnect_0_oil_temp_s1_chipselect),                     //                                           .chipselect
		.sysid_c001_control_slave_address                 (mm_interconnect_0_sysid_c001_control_slave_address),           //                   sysid_c001_control_slave.address
		.sysid_c001_control_slave_readdata                (mm_interconnect_0_sysid_c001_control_slave_readdata),          //                                           .readdata
		.wrn_s1_address                                   (mm_interconnect_0_wrn_s1_address),                             //                                     wrn_s1.address
		.wrn_s1_write                                     (mm_interconnect_0_wrn_s1_write),                               //                                           .write
		.wrn_s1_readdata                                  (mm_interconnect_0_wrn_s1_readdata),                            //                                           .readdata
		.wrn_s1_writedata                                 (mm_interconnect_0_wrn_s1_writedata),                           //                                           .writedata
		.wrn_s1_chipselect                                (mm_interconnect_0_wrn_s1_chipselect)                           //                                           .chipselect
	);

	controller_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_qsys_0_d_irq_irq)          //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in0.reset
		.reset_in1      (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),             // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),         //          .reset_req
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_in2      (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

endmodule
