// controller_tb.v

// Generated using ACDS version 13.1 162 at 2018.07.24.21:25:12

`timescale 1 ps / 1 ps
module controller_tb (
	);

	wire         controller_inst_clock_50_bfm_clk_clk;                    // controller_inst_clock_50_bfm:clk -> [controller_inst:clock_50_clk, controller_inst_reset_bfm:clk]
	wire         controller_inst_reset_bfm_reset_reset;                   // controller_inst_reset_bfm:reset -> controller_inst:reset_reset_n
	wire   [0:0] controller_inst_daylight_bfm_conduit_export;             // controller_inst_daylight_bfm:sig_export -> controller_inst:daylight_export
	wire  [31:0] controller_inst_tc1_m_export;                            // controller_inst:tc1_m_export -> controller_inst_tc1_m_bfm:sig_export
	wire  [31:0] controller_inst_tc2_m_export;                            // controller_inst:tc2_m_export -> controller_inst_tc2_m_bfm:sig_export
	wire  [31:0] controller_inst_tc3_m_export;                            // controller_inst:tc3_m_export -> controller_inst_tc3_m_bfm:sig_export
	wire  [31:0] controller_inst_tc4_m_export;                            // controller_inst:tc4_m_export -> controller_inst_tc4_m_bfm:sig_export
	wire   [3:0] controller_inst_tc_reset_export;                         // controller_inst:tc_reset_export -> controller_inst_tc_reset_bfm:sig_export
	wire  [24:0] controller_inst_tc1_status_bfm_conduit_export;           // controller_inst_tc1_status_bfm:sig_export -> controller_inst:tc1_status_export
	wire  [24:0] controller_inst_tc2_status_bfm_conduit_export;           // controller_inst_tc2_status_bfm:sig_export -> controller_inst:tc2_status_export
	wire  [24:0] controller_inst_tc3_status_bfm_conduit_export;           // controller_inst_tc3_status_bfm:sig_export -> controller_inst:tc3_status_export
	wire  [24:0] controller_inst_tc4_status_bfm_conduit_export;           // controller_inst_tc4_status_bfm:sig_export -> controller_inst:tc4_status_export
	wire   [7:0] controller_inst_uart1_w_data_export;                     // controller_inst:uart1_w_data_export -> controller_inst_uart1_w_data_bfm:sig_export
	wire   [2:0] controller_inst_uart1_reset_control_export;              // controller_inst:uart1_reset_control_export -> controller_inst_uart1_reset_control_bfm:sig_export
	wire   [1:0] controller_inst_uart1_wr_control_export;                 // controller_inst:uart1_wr_control_export -> controller_inst_uart1_wr_control_bfm:sig_export
	wire  [21:0] controller_inst_uart1_baud_control_export;               // controller_inst:uart1_baud_control_export -> controller_inst_uart1_baud_control_bfm:sig_export
	wire   [7:0] controller_inst_uart1_r_data_bfm_conduit_export;         // controller_inst_uart1_r_data_bfm:sig_export -> controller_inst:uart1_r_data_export
	wire   [7:0] controller_inst_uart1_rx_counter_bfm_conduit_export;     // controller_inst_uart1_rx_counter_bfm:sig_export -> controller_inst:uart1_rx_counter_export
	wire   [2:0] controller_inst_uart1_tx_counter_bfm_conduit_export;     // controller_inst_uart1_tx_counter_bfm:sig_export -> controller_inst:uart1_tx_counter_export
	wire   [7:0] controller_inst_uart1_status_control_bfm_conduit_export; // controller_inst_uart1_status_control_bfm:sig_export -> controller_inst:uart1_status_control_export
	wire  [13:0] controller_inst_bcd1_bin_export;                         // controller_inst:bcd1_bin_export -> controller_inst_bcd1_bin_bfm:sig_export
	wire   [2:0] controller_inst_bcd1_control_export;                     // controller_inst:bcd1_control_export -> controller_inst_bcd1_control_bfm:sig_export
	wire  [15:0] controller_inst_bcd1_bcd_bfm_conduit_export;             // controller_inst_bcd1_bcd_bfm:sig_export -> controller_inst:bcd1_bcd_export
	wire   [7:0] controller_inst_bcd1_counter_bfm_conduit_export;         // controller_inst_bcd1_counter_bfm:sig_export -> controller_inst:bcd1_counter_export
	wire   [1:0] controller_inst_bcd1_status_bfm_conduit_export;          // controller_inst_bcd1_status_bfm:sig_export -> controller_inst:bcd1_status_export
	wire   [7:0] controller_inst_warn_pwm_brightness_export;              // controller_inst:warn_pwm_brightness_export -> controller_inst_warn_pwm_brightness_bfm:sig_export
	wire   [3:0] controller_inst_status_led_en_export;                    // controller_inst:status_led_en_export -> controller_inst_status_led_en_bfm:sig_export
	wire   [1:0] controller_inst_warn_pwm_control_export;                 // controller_inst:warn_pwm_control_export -> controller_inst_warn_pwm_control_bfm:sig_export
	wire   [7:0] controller_inst_sseg_brightness_boost_export;            // controller_inst:sseg_brightness_boost_export -> controller_inst_sseg_brightness_boost_bfm:sig_export
	wire   [7:0] controller_inst_sseg_brightness_afr_export;              // controller_inst:sseg_brightness_afr_export -> controller_inst_sseg_brightness_afr_bfm:sig_export
	wire   [7:0] controller_inst_sseg_brightness_oil_export;              // controller_inst:sseg_brightness_oil_export -> controller_inst_sseg_brightness_oil_bfm:sig_export
	wire   [7:0] controller_inst_sseg_brightness_coolant_export;          // controller_inst:sseg_brightness_coolant_export -> controller_inst_sseg_brightness_coolant_bfm:sig_export
	wire   [1:0] controller_inst_sseg_sel_addr_export;                    // controller_inst:sseg_sel_addr_export -> controller_inst_sseg_sel_addr_bfm:sig_export
	wire   [4:0] controller_inst_sseg_reset_control_export;               // controller_inst:sseg_reset_control_export -> controller_inst_sseg_reset_control_bfm:sig_export
	wire   [3:0] controller_inst_sseg_wr_control_export;                  // controller_inst:sseg_wr_control_export -> controller_inst_sseg_wr_control_bfm:sig_export
	wire   [6:0] controller_inst_sseg_wr_val_export;                      // controller_inst:sseg_wr_val_export -> controller_inst_sseg_wr_val_bfm:sig_export
	wire   [7:0] controller_inst_sseg_counter_bfm_conduit_export;         // controller_inst_sseg_counter_bfm:sig_export -> controller_inst:sseg_counter_export
	wire   [0:0] controller_inst_sseg_counter_of_bfm_conduit_export;      // controller_inst_sseg_counter_of_bfm:sig_export -> controller_inst:sseg_counter_of_export
	wire   [7:0] controller_inst_leds_boost_brightness_export;            // controller_inst:leds_boost_brightness_export -> controller_inst_leds_boost_brightness_bfm:sig_export
	wire   [7:0] controller_inst_leds_afr_brightness_export;              // controller_inst:leds_afr_brightness_export -> controller_inst_leds_afr_brightness_bfm:sig_export
	wire   [5:0] controller_inst_leds_afr_sel_addr_export;                // controller_inst:leds_afr_sel_addr_export -> controller_inst_leds_afr_sel_addr_bfm:sig_export
	wire   [5:0] controller_inst_leds_boost_sel_addr_export;              // controller_inst:leds_boost_sel_addr_export -> controller_inst_leds_boost_sel_addr_bfm:sig_export
	wire   [3:0] controller_inst_leds_reset_control_export;               // controller_inst:leds_reset_control_export -> controller_inst_leds_reset_control_bfm:sig_export
	wire   [1:0] controller_inst_leds_afr_control_export;                 // controller_inst:leds_afr_control_export -> controller_inst_leds_afr_control_bfm:sig_export
	wire   [7:0] controller_inst_leds_boost_counter_bfm_conduit_export;   // controller_inst_leds_boost_counter_bfm:sig_export -> controller_inst:leds_boost_counter_export
	wire   [1:0] controller_inst_leds_boost_control_export;               // controller_inst:leds_boost_control_export -> controller_inst_leds_boost_control_bfm:sig_export
	wire   [7:0] controller_inst_leds_afr_counter_bfm_conduit_export;     // controller_inst_leds_afr_counter_bfm:sig_export -> controller_inst:leds_afr_counter_export
	wire   [1:0] controller_inst_leds_counter_status_bfm_conduit_export;  // controller_inst_leds_counter_status_bfm:sig_export -> controller_inst:leds_counter_status_export
	wire  [15:0] controller_inst_uart1_dvsr_export;                       // controller_inst:uart1_dvsr_export -> controller_inst_uart1_dvsr_bfm:sig_export

	controller controller_inst (
		.clock_50_clk                   (controller_inst_clock_50_bfm_clk_clk),                    //                clock_50.clk
		.daylight_export                (controller_inst_daylight_bfm_conduit_export),             //                daylight.export
		.tc1_m_export                   (controller_inst_tc1_m_export),                            //                   tc1_m.export
		.tc2_m_export                   (controller_inst_tc2_m_export),                            //                   tc2_m.export
		.tc3_m_export                   (controller_inst_tc3_m_export),                            //                   tc3_m.export
		.tc4_m_export                   (controller_inst_tc4_m_export),                            //                   tc4_m.export
		.tc_reset_export                (controller_inst_tc_reset_export),                         //                tc_reset.export
		.tc1_status_export              (controller_inst_tc1_status_bfm_conduit_export),           //              tc1_status.export
		.tc2_status_export              (controller_inst_tc2_status_bfm_conduit_export),           //              tc2_status.export
		.tc3_status_export              (controller_inst_tc3_status_bfm_conduit_export),           //              tc3_status.export
		.tc4_status_export              (controller_inst_tc4_status_bfm_conduit_export),           //              tc4_status.export
		.uart1_w_data_export            (controller_inst_uart1_w_data_export),                     //            uart1_w_data.export
		.uart1_reset_control_export     (controller_inst_uart1_reset_control_export),              //     uart1_reset_control.export
		.uart1_wr_control_export        (controller_inst_uart1_wr_control_export),                 //        uart1_wr_control.export
		.uart1_baud_control_export      (controller_inst_uart1_baud_control_export),               //      uart1_baud_control.export
		.uart1_r_data_export            (controller_inst_uart1_r_data_bfm_conduit_export),         //            uart1_r_data.export
		.uart1_rx_counter_export        (controller_inst_uart1_rx_counter_bfm_conduit_export),     //        uart1_rx_counter.export
		.uart1_tx_counter_export        (controller_inst_uart1_tx_counter_bfm_conduit_export),     //        uart1_tx_counter.export
		.uart1_status_control_export    (controller_inst_uart1_status_control_bfm_conduit_export), //    uart1_status_control.export
		.bcd1_bin_export                (controller_inst_bcd1_bin_export),                         //                bcd1_bin.export
		.bcd1_control_export            (controller_inst_bcd1_control_export),                     //            bcd1_control.export
		.bcd1_bcd_export                (controller_inst_bcd1_bcd_bfm_conduit_export),             //                bcd1_bcd.export
		.bcd1_counter_export            (controller_inst_bcd1_counter_bfm_conduit_export),         //            bcd1_counter.export
		.bcd1_status_export             (controller_inst_bcd1_status_bfm_conduit_export),          //             bcd1_status.export
		.warn_pwm_brightness_export     (controller_inst_warn_pwm_brightness_export),              //     warn_pwm_brightness.export
		.status_led_en_export           (controller_inst_status_led_en_export),                    //           status_led_en.export
		.warn_pwm_control_export        (controller_inst_warn_pwm_control_export),                 //        warn_pwm_control.export
		.sseg_brightness_boost_export   (controller_inst_sseg_brightness_boost_export),            //   sseg_brightness_boost.export
		.sseg_brightness_afr_export     (controller_inst_sseg_brightness_afr_export),              //     sseg_brightness_afr.export
		.sseg_brightness_oil_export     (controller_inst_sseg_brightness_oil_export),              //     sseg_brightness_oil.export
		.sseg_brightness_coolant_export (controller_inst_sseg_brightness_coolant_export),          // sseg_brightness_coolant.export
		.sseg_sel_addr_export           (controller_inst_sseg_sel_addr_export),                    //           sseg_sel_addr.export
		.sseg_reset_control_export      (controller_inst_sseg_reset_control_export),               //      sseg_reset_control.export
		.sseg_wr_control_export         (controller_inst_sseg_wr_control_export),                  //         sseg_wr_control.export
		.sseg_wr_val_export             (controller_inst_sseg_wr_val_export),                      //             sseg_wr_val.export
		.sseg_counter_export            (controller_inst_sseg_counter_bfm_conduit_export),         //            sseg_counter.export
		.sseg_counter_of_export         (controller_inst_sseg_counter_of_bfm_conduit_export),      //         sseg_counter_of.export
		.leds_boost_brightness_export   (controller_inst_leds_boost_brightness_export),            //   leds_boost_brightness.export
		.leds_afr_brightness_export     (controller_inst_leds_afr_brightness_export),              //     leds_afr_brightness.export
		.leds_afr_sel_addr_export       (controller_inst_leds_afr_sel_addr_export),                //       leds_afr_sel_addr.export
		.leds_boost_sel_addr_export     (controller_inst_leds_boost_sel_addr_export),              //     leds_boost_sel_addr.export
		.leds_reset_control_export      (controller_inst_leds_reset_control_export),               //      leds_reset_control.export
		.leds_afr_control_export        (controller_inst_leds_afr_control_export),                 //        leds_afr_control.export
		.leds_boost_counter_export      (controller_inst_leds_boost_counter_bfm_conduit_export),   //      leds_boost_counter.export
		.leds_boost_control_export      (controller_inst_leds_boost_control_export),               //      leds_boost_control.export
		.leds_afr_counter_export        (controller_inst_leds_afr_counter_bfm_conduit_export),     //        leds_afr_counter.export
		.leds_counter_status_export     (controller_inst_leds_counter_status_bfm_conduit_export),  //     leds_counter_status.export
		.reset_reset_n                  (controller_inst_reset_bfm_reset_reset),                   //                   reset.reset_n
		.uart1_dvsr_export              (controller_inst_uart1_dvsr_export)                        //              uart1_dvsr.export
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) controller_inst_clock_50_bfm (
		.clk (controller_inst_clock_50_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) controller_inst_reset_bfm (
		.reset (controller_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (controller_inst_clock_50_bfm_clk_clk)   //   clk.clk
	);

	altera_conduit_bfm controller_inst_daylight_bfm (
		.sig_export (controller_inst_daylight_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0002 controller_inst_tc1_m_bfm (
		.sig_export (controller_inst_tc1_m_export)  // conduit.export
	);

	altera_conduit_bfm_0002 controller_inst_tc2_m_bfm (
		.sig_export (controller_inst_tc2_m_export)  // conduit.export
	);

	altera_conduit_bfm_0002 controller_inst_tc3_m_bfm (
		.sig_export (controller_inst_tc3_m_export)  // conduit.export
	);

	altera_conduit_bfm_0002 controller_inst_tc4_m_bfm (
		.sig_export (controller_inst_tc4_m_export)  // conduit.export
	);

	altera_conduit_bfm_0003 controller_inst_tc_reset_bfm (
		.sig_export (controller_inst_tc_reset_export)  // conduit.export
	);

	altera_conduit_bfm_0004 controller_inst_tc1_status_bfm (
		.sig_export (controller_inst_tc1_status_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0004 controller_inst_tc2_status_bfm (
		.sig_export (controller_inst_tc2_status_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0004 controller_inst_tc3_status_bfm (
		.sig_export (controller_inst_tc3_status_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0004 controller_inst_tc4_status_bfm (
		.sig_export (controller_inst_tc4_status_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0005 controller_inst_uart1_w_data_bfm (
		.sig_export (controller_inst_uart1_w_data_export)  // conduit.export
	);

	altera_conduit_bfm_0006 controller_inst_uart1_reset_control_bfm (
		.sig_export (controller_inst_uart1_reset_control_export)  // conduit.export
	);

	altera_conduit_bfm_0007 controller_inst_uart1_wr_control_bfm (
		.sig_export (controller_inst_uart1_wr_control_export)  // conduit.export
	);

	altera_conduit_bfm_0008 controller_inst_uart1_baud_control_bfm (
		.sig_export (controller_inst_uart1_baud_control_export)  // conduit.export
	);

	altera_conduit_bfm_0009 controller_inst_uart1_r_data_bfm (
		.sig_export (controller_inst_uart1_r_data_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0009 controller_inst_uart1_rx_counter_bfm (
		.sig_export (controller_inst_uart1_rx_counter_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0010 controller_inst_uart1_tx_counter_bfm (
		.sig_export (controller_inst_uart1_tx_counter_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0009 controller_inst_uart1_status_control_bfm (
		.sig_export (controller_inst_uart1_status_control_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0011 controller_inst_bcd1_bin_bfm (
		.sig_export (controller_inst_bcd1_bin_export)  // conduit.export
	);

	altera_conduit_bfm_0006 controller_inst_bcd1_control_bfm (
		.sig_export (controller_inst_bcd1_control_export)  // conduit.export
	);

	altera_conduit_bfm_0012 controller_inst_bcd1_bcd_bfm (
		.sig_export (controller_inst_bcd1_bcd_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0009 controller_inst_bcd1_counter_bfm (
		.sig_export (controller_inst_bcd1_counter_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0013 controller_inst_bcd1_status_bfm (
		.sig_export (controller_inst_bcd1_status_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0005 controller_inst_warn_pwm_brightness_bfm (
		.sig_export (controller_inst_warn_pwm_brightness_export)  // conduit.export
	);

	altera_conduit_bfm_0003 controller_inst_status_led_en_bfm (
		.sig_export (controller_inst_status_led_en_export)  // conduit.export
	);

	altera_conduit_bfm_0007 controller_inst_warn_pwm_control_bfm (
		.sig_export (controller_inst_warn_pwm_control_export)  // conduit.export
	);

	altera_conduit_bfm_0005 controller_inst_sseg_brightness_boost_bfm (
		.sig_export (controller_inst_sseg_brightness_boost_export)  // conduit.export
	);

	altera_conduit_bfm_0005 controller_inst_sseg_brightness_afr_bfm (
		.sig_export (controller_inst_sseg_brightness_afr_export)  // conduit.export
	);

	altera_conduit_bfm_0005 controller_inst_sseg_brightness_oil_bfm (
		.sig_export (controller_inst_sseg_brightness_oil_export)  // conduit.export
	);

	altera_conduit_bfm_0005 controller_inst_sseg_brightness_coolant_bfm (
		.sig_export (controller_inst_sseg_brightness_coolant_export)  // conduit.export
	);

	altera_conduit_bfm_0007 controller_inst_sseg_sel_addr_bfm (
		.sig_export (controller_inst_sseg_sel_addr_export)  // conduit.export
	);

	altera_conduit_bfm_0014 controller_inst_sseg_reset_control_bfm (
		.sig_export (controller_inst_sseg_reset_control_export)  // conduit.export
	);

	altera_conduit_bfm_0003 controller_inst_sseg_wr_control_bfm (
		.sig_export (controller_inst_sseg_wr_control_export)  // conduit.export
	);

	altera_conduit_bfm_0015 controller_inst_sseg_wr_val_bfm (
		.sig_export (controller_inst_sseg_wr_val_export)  // conduit.export
	);

	altera_conduit_bfm_0009 controller_inst_sseg_counter_bfm (
		.sig_export (controller_inst_sseg_counter_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm controller_inst_sseg_counter_of_bfm (
		.sig_export (controller_inst_sseg_counter_of_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0005 controller_inst_leds_boost_brightness_bfm (
		.sig_export (controller_inst_leds_boost_brightness_export)  // conduit.export
	);

	altera_conduit_bfm_0005 controller_inst_leds_afr_brightness_bfm (
		.sig_export (controller_inst_leds_afr_brightness_export)  // conduit.export
	);

	altera_conduit_bfm_0016 controller_inst_leds_afr_sel_addr_bfm (
		.sig_export (controller_inst_leds_afr_sel_addr_export)  // conduit.export
	);

	altera_conduit_bfm_0016 controller_inst_leds_boost_sel_addr_bfm (
		.sig_export (controller_inst_leds_boost_sel_addr_export)  // conduit.export
	);

	altera_conduit_bfm_0003 controller_inst_leds_reset_control_bfm (
		.sig_export (controller_inst_leds_reset_control_export)  // conduit.export
	);

	altera_conduit_bfm_0007 controller_inst_leds_afr_control_bfm (
		.sig_export (controller_inst_leds_afr_control_export)  // conduit.export
	);

	altera_conduit_bfm_0009 controller_inst_leds_boost_counter_bfm (
		.sig_export (controller_inst_leds_boost_counter_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0007 controller_inst_leds_boost_control_bfm (
		.sig_export (controller_inst_leds_boost_control_export)  // conduit.export
	);

	altera_conduit_bfm_0009 controller_inst_leds_afr_counter_bfm (
		.sig_export (controller_inst_leds_afr_counter_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0013 controller_inst_leds_counter_status_bfm (
		.sig_export (controller_inst_leds_counter_status_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0017 controller_inst_uart1_dvsr_bfm (
		.sig_export (controller_inst_uart1_dvsr_export)  // conduit.export
	);

endmodule
