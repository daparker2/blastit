// controller_tb.v

// Generated using ACDS version 13.1 162 at 2018.07.17.20:32:36

`timescale 1 ps / 1 ps
module controller_tb (
	);

	wire        controller_inst_clock_50_bfm_clk_clk;  // controller_inst_clock_50_bfm:clk -> [controller_inst:clock_50_clk, controller_inst_reset_bfm:clk]
	wire        controller_inst_reset_bfm_reset_reset; // controller_inst_reset_bfm:reset -> controller_inst:reset_reset_n
	wire  [2:0] controller_inst_warning_en_export;     // controller_inst:warning_en_export -> controller_inst_warning_en_bfm:sig_export

	controller controller_inst (
		.clock_50_clk      (controller_inst_clock_50_bfm_clk_clk),  //   clock_50.clk
		.warning_en_export (controller_inst_warning_en_export),     // warning_en.export
		.reset_reset_n     (controller_inst_reset_bfm_reset_reset)  //      reset.reset_n
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) controller_inst_clock_50_bfm (
		.clk (controller_inst_clock_50_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) controller_inst_reset_bfm (
		.reset (controller_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (controller_inst_clock_50_bfm_clk_clk)   //   clk.clk
	);

	altera_conduit_bfm controller_inst_warning_en_bfm (
		.sig_export (controller_inst_warning_en_export)  // conduit.export
	);

endmodule
