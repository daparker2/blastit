module sseg
(
	input wire[3:0] num,
	output reg[6:0] hex
);

	always @*
	begin
		case (num)
			4'h0: hex[6:0] = 7'b1000000;
			4'h1: hex[6:0] = 7'b1111001;
			4'h2: hex[6:0] = 7'b0100100;
			4'h3: hex[6:0] = 7'b0110000;
			4'h4: hex[6:0] = 7'b0011001;
			4'h5: hex[6:0] = 7'b0010010;
			4'h6: hex[6:0] = 7'b0000010;
			4'h7: hex[6:0] = 7'b1111000;
			4'h8: hex[6:0] = 7'b0000000;
			4'h9: hex[6:0] = 7'b0010000;
			4'ha: hex[6:0] = 7'b0001000;
			4'hb: hex[6:0] = 7'b0000011;
			4'hc: hex[6:0] = 7'b0100111;
			4'hd: hex[6:0] = 7'b0100001;
			4'he: hex[6:0] = 7'b0000110;
			4'hf: hex[6:0] = 7'b0001110;
			default: hex[6:0] = 7'b0101100;
		endcase
	end

endmodule