// controller_tb.v

// Generated using ACDS version 13.1 162 at 2018.10.06.18:06:30

`timescale 1 ps / 1 ps
module controller_tb (
	);

	wire    controller_inst_clock_50_bfm_clk_clk;  // controller_inst_clock_50_bfm:clk -> [controller_inst:clock_50_clk, controller_inst_reset_bfm:clk]
	wire    controller_inst_reset_bfm_reset_reset; // controller_inst_reset_bfm:reset -> controller_inst:reset_reset_n

	controller controller_inst (
		.clock_50_clk                (controller_inst_clock_50_bfm_clk_clk),  //             clock_50.clk
		.daylight_export             (),                                      //             daylight.export
		.tc1_m_export                (),                                      //                tc1_m.export
		.tc2_m_export                (),                                      //                tc2_m.export
		.tc3_m_export                (),                                      //                tc3_m.export
		.tc4_m_export                (),                                      //                tc4_m.export
		.tc_reset_control_export     (),                                      //     tc_reset_control.export
		.tc1_status_export           (),                                      //           tc1_status.export
		.tc2_status_export           (),                                      //           tc2_status.export
		.tc3_status_export           (),                                      //           tc3_status.export
		.tc4_status_export           (),                                      //           tc4_status.export
		.uart1_w_data_export         (),                                      //         uart1_w_data.export
		.uart1_reset_control_export  (),                                      //  uart1_reset_control.export
		.uart1_wr_control_export     (),                                      //     uart1_wr_control.export
		.uart1_baud_control_export   (),                                      //   uart1_baud_control.export
		.uart1_r_data_export         (),                                      //         uart1_r_data.export
		.uart1_rx_counter_export     (),                                      //     uart1_rx_counter.export
		.uart1_tx_counter_export     (),                                      //     uart1_tx_counter.export
		.uart1_status_control_export (),                                      // uart1_status_control.export
		.bcd1_bin_export             (),                                      //             bcd1_bin.export
		.bcd1_control_export         (),                                      //         bcd1_control.export
		.bcd1_bcd_export             (),                                      //             bcd1_bcd.export
		.bcd1_counter_export         (),                                      //         bcd1_counter.export
		.bcd1_status_export          (),                                      //          bcd1_status.export
		.warn_pwm_brightness_export  (),                                      //  warn_pwm_brightness.export
		.status_led_en_export        (),                                      //        status_led_en.export
		.warn_pwm_control_export     (),                                      //     warn_pwm_control.export
		.sseg_brightness_export      (),                                      //      sseg_brightness.export
		.sseg_reset_control_export   (),                                      //   sseg_reset_control.export
		.sseg_wr_val_export          (),                                      //          sseg_wr_val.export
		.sseg_counter_export         (),                                      //         sseg_counter.export
		.sseg_counter_of_export      (),                                      //      sseg_counter_of.export
		.leds1_brightness_export     (),                                      //     leds1_brightness.export
		.leds1_wr_val_export         (),                                      //         leds1_wr_val.export
		.leds1_counter_export        (),                                      //        leds1_counter.export
		.leds1_reset_control_export  (),                                      //  leds1_reset_control.export
		.leds1_counter_of_export     (),                                      //     leds1_counter_of.export
		.reset_reset_n               (controller_inst_reset_bfm_reset_reset), //                reset.reset_n
		.uart1_dvsr_export           (),                                      //           uart1_dvsr.export
		.rc1_control_export          (),                                      //          rc1_control.export
		.rc1_ready_export            (),                                      //            rc1_ready.export
		.led_period_export           (),                                      //           led_period.export
		.leds2_reset_control_export  (),                                      //  leds2_reset_control.export
		.leds2_wr_val_export         (),                                      //         leds2_wr_val.export
		.leds2_counter_export        (),                                      //        leds2_counter.export
		.leds2_counter_of_export     (),                                      //     leds2_counter_of.export
		.leds2_brightness_export     ()                                       //     leds2_brightness.export
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) controller_inst_clock_50_bfm (
		.clk (controller_inst_clock_50_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) controller_inst_reset_bfm (
		.reset (controller_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (controller_inst_clock_50_bfm_clk_clk)   //   clk.clk
	);

endmodule
