// controller.v

// Generated using ACDS version 13.1 162 at 2018.09.21.22:23:51

`timescale 1 ps / 1 ps
module controller (
		input  wire        clock_50_clk,                //             clock_50.clk
		input  wire        daylight_export,             //             daylight.export
		output wire [31:0] tc1_m_export,                //                tc1_m.export
		output wire [31:0] tc2_m_export,                //                tc2_m.export
		output wire [31:0] tc3_m_export,                //                tc3_m.export
		output wire [31:0] tc4_m_export,                //                tc4_m.export
		output wire [3:0]  tc_reset_control_export,     //     tc_reset_control.export
		input  wire [24:0] tc1_status_export,           //           tc1_status.export
		input  wire [24:0] tc2_status_export,           //           tc2_status.export
		input  wire [24:0] tc3_status_export,           //           tc3_status.export
		input  wire [24:0] tc4_status_export,           //           tc4_status.export
		output wire [7:0]  uart1_w_data_export,         //         uart1_w_data.export
		output wire [2:0]  uart1_reset_control_export,  //  uart1_reset_control.export
		output wire [1:0]  uart1_wr_control_export,     //     uart1_wr_control.export
		output wire [21:0] uart1_baud_control_export,   //   uart1_baud_control.export
		input  wire [7:0]  uart1_r_data_export,         //         uart1_r_data.export
		input  wire [7:0]  uart1_rx_counter_export,     //     uart1_rx_counter.export
		input  wire [7:0]  uart1_tx_counter_export,     //     uart1_tx_counter.export
		input  wire [9:0]  uart1_status_control_export, // uart1_status_control.export
		output wire [14:0] bcd1_bin_export,             //             bcd1_bin.export
		output wire [2:0]  bcd1_control_export,         //         bcd1_control.export
		input  wire [15:0] bcd1_bcd_export,             //             bcd1_bcd.export
		input  wire [7:0]  bcd1_counter_export,         //         bcd1_counter.export
		input  wire [1:0]  bcd1_status_export,          //          bcd1_status.export
		output wire [7:0]  warn_pwm_brightness_export,  //  warn_pwm_brightness.export
		output wire [3:0]  status_led_en_export,        //        status_led_en.export
		output wire [1:0]  warn_pwm_control_export,     //     warn_pwm_control.export
		output wire [7:0]  sseg_brightness_export,      //      sseg_brightness.export
		output wire [1:0]  sseg_reset_control_export,   //   sseg_reset_control.export
		output wire [12:0] sseg_wr_val_export,          //          sseg_wr_val.export
		input  wire [7:0]  sseg_counter_export,         //         sseg_counter.export
		input  wire        sseg_counter_of_export,      //      sseg_counter_of.export
		output wire [7:0]  leds1_brightness_export,     //     leds1_brightness.export
		output wire [9:0]  leds1_wr_val_export,         //         leds1_wr_val.export
		input  wire [7:0]  leds1_counter_export,        //        leds1_counter.export
		output wire [1:0]  leds1_reset_control_export,  //  leds1_reset_control.export
		input  wire        leds1_counter_of_export,     //     leds1_counter_of.export
		input  wire        reset_reset_n,               //                reset.reset_n
		output wire [15:0] uart1_dvsr_export,           //           uart1_dvsr.export
		output wire [24:0] rc1_control_export,          //          rc1_control.export
		input  wire        rc1_ready_export,            //            rc1_ready.export
		output wire [23:0] led_period_export,           //           led_period.export
		output wire [1:0]  leds2_reset_control_export,  //  leds2_reset_control.export
		output wire [9:0]  leds2_wr_val_export,         //         leds2_wr_val.export
		input  wire [7:0]  leds2_counter_export,        //        leds2_counter.export
		input  wire        leds2_counter_of_export,     //     leds2_counter_of.export
		output wire [7:0]  leds2_brightness_export      //     leds2_brightness.export
	);

	wire  [31:0] mm_interconnect_0_tc3_m_s1_writedata;                        // mm_interconnect_0:tc3_m_s1_writedata -> tc3_m:writedata
	wire   [1:0] mm_interconnect_0_tc3_m_s1_address;                          // mm_interconnect_0:tc3_m_s1_address -> tc3_m:address
	wire         mm_interconnect_0_tc3_m_s1_chipselect;                       // mm_interconnect_0:tc3_m_s1_chipselect -> tc3_m:chipselect
	wire         mm_interconnect_0_tc3_m_s1_write;                            // mm_interconnect_0:tc3_m_s1_write -> tc3_m:write_n
	wire  [31:0] mm_interconnect_0_tc3_m_s1_readdata;                         // tc3_m:readdata -> mm_interconnect_0:tc3_m_s1_readdata
	wire  [31:0] mm_interconnect_0_leds1_reset_control_s1_writedata;          // mm_interconnect_0:leds1_reset_control_s1_writedata -> leds1_reset_control:writedata
	wire   [1:0] mm_interconnect_0_leds1_reset_control_s1_address;            // mm_interconnect_0:leds1_reset_control_s1_address -> leds1_reset_control:address
	wire         mm_interconnect_0_leds1_reset_control_s1_chipselect;         // mm_interconnect_0:leds1_reset_control_s1_chipselect -> leds1_reset_control:chipselect
	wire         mm_interconnect_0_leds1_reset_control_s1_write;              // mm_interconnect_0:leds1_reset_control_s1_write -> leds1_reset_control:write_n
	wire  [31:0] mm_interconnect_0_leds1_reset_control_s1_readdata;           // leds1_reset_control:readdata -> mm_interconnect_0:leds1_reset_control_s1_readdata
	wire  [31:0] mm_interconnect_0_tc_reset_control_s1_writedata;             // mm_interconnect_0:tc_reset_control_s1_writedata -> tc_reset_control:writedata
	wire   [1:0] mm_interconnect_0_tc_reset_control_s1_address;               // mm_interconnect_0:tc_reset_control_s1_address -> tc_reset_control:address
	wire         mm_interconnect_0_tc_reset_control_s1_chipselect;            // mm_interconnect_0:tc_reset_control_s1_chipselect -> tc_reset_control:chipselect
	wire         mm_interconnect_0_tc_reset_control_s1_write;                 // mm_interconnect_0:tc_reset_control_s1_write -> tc_reset_control:write_n
	wire  [31:0] mm_interconnect_0_tc_reset_control_s1_readdata;              // tc_reset_control:readdata -> mm_interconnect_0:tc_reset_control_s1_readdata
	wire   [1:0] mm_interconnect_0_leds2_counter_s1_address;                  // mm_interconnect_0:leds2_counter_s1_address -> leds2_counter:address
	wire  [31:0] mm_interconnect_0_leds2_counter_s1_readdata;                 // leds2_counter:readdata -> mm_interconnect_0:leds2_counter_s1_readdata
	wire  [31:0] mm_interconnect_0_tc4_m_s1_writedata;                        // mm_interconnect_0:tc4_m_s1_writedata -> tc4_m:writedata
	wire   [1:0] mm_interconnect_0_tc4_m_s1_address;                          // mm_interconnect_0:tc4_m_s1_address -> tc4_m:address
	wire         mm_interconnect_0_tc4_m_s1_chipselect;                       // mm_interconnect_0:tc4_m_s1_chipselect -> tc4_m:chipselect
	wire         mm_interconnect_0_tc4_m_s1_write;                            // mm_interconnect_0:tc4_m_s1_write -> tc4_m:write_n
	wire  [31:0] mm_interconnect_0_tc4_m_s1_readdata;                         // tc4_m:readdata -> mm_interconnect_0:tc4_m_s1_readdata
	wire   [1:0] mm_interconnect_0_tc1_status_s1_address;                     // mm_interconnect_0:tc1_status_s1_address -> tc1_status:address
	wire  [31:0] mm_interconnect_0_tc1_status_s1_readdata;                    // tc1_status:readdata -> mm_interconnect_0:tc1_status_s1_readdata
	wire   [1:0] mm_interconnect_0_uart1_status_control_s1_address;           // mm_interconnect_0:uart1_status_control_s1_address -> uart1_status_control:address
	wire  [31:0] mm_interconnect_0_uart1_status_control_s1_readdata;          // uart1_status_control:readdata -> mm_interconnect_0:uart1_status_control_s1_readdata
	wire   [1:0] mm_interconnect_0_tc4_status_s1_address;                     // mm_interconnect_0:tc4_status_s1_address -> tc4_status:address
	wire  [31:0] mm_interconnect_0_tc4_status_s1_readdata;                    // tc4_status:readdata -> mm_interconnect_0:tc4_status_s1_readdata
	wire  [31:0] mm_interconnect_0_rc1_control_s1_writedata;                  // mm_interconnect_0:rc1_control_s1_writedata -> rc1_control:writedata
	wire   [1:0] mm_interconnect_0_rc1_control_s1_address;                    // mm_interconnect_0:rc1_control_s1_address -> rc1_control:address
	wire         mm_interconnect_0_rc1_control_s1_chipselect;                 // mm_interconnect_0:rc1_control_s1_chipselect -> rc1_control:chipselect
	wire         mm_interconnect_0_rc1_control_s1_write;                      // mm_interconnect_0:rc1_control_s1_write -> rc1_control:write_n
	wire  [31:0] mm_interconnect_0_rc1_control_s1_readdata;                   // rc1_control:readdata -> mm_interconnect_0:rc1_control_s1_readdata
	wire   [1:0] mm_interconnect_0_uart1_rx_counter_s1_address;               // mm_interconnect_0:uart1_rx_counter_s1_address -> uart1_rx_counter:address
	wire  [31:0] mm_interconnect_0_uart1_rx_counter_s1_readdata;              // uart1_rx_counter:readdata -> mm_interconnect_0:uart1_rx_counter_s1_readdata
	wire  [31:0] mm_interconnect_0_uart1_w_data_s1_writedata;                 // mm_interconnect_0:uart1_w_data_s1_writedata -> uart1_w_data:writedata
	wire   [1:0] mm_interconnect_0_uart1_w_data_s1_address;                   // mm_interconnect_0:uart1_w_data_s1_address -> uart1_w_data:address
	wire         mm_interconnect_0_uart1_w_data_s1_chipselect;                // mm_interconnect_0:uart1_w_data_s1_chipselect -> uart1_w_data:chipselect
	wire         mm_interconnect_0_uart1_w_data_s1_write;                     // mm_interconnect_0:uart1_w_data_s1_write -> uart1_w_data:write_n
	wire  [31:0] mm_interconnect_0_uart1_w_data_s1_readdata;                  // uart1_w_data:readdata -> mm_interconnect_0:uart1_w_data_s1_readdata
	wire  [31:0] mm_interconnect_0_uart1_wr_control_s1_writedata;             // mm_interconnect_0:uart1_wr_control_s1_writedata -> uart1_wr_control:writedata
	wire   [1:0] mm_interconnect_0_uart1_wr_control_s1_address;               // mm_interconnect_0:uart1_wr_control_s1_address -> uart1_wr_control:address
	wire         mm_interconnect_0_uart1_wr_control_s1_chipselect;            // mm_interconnect_0:uart1_wr_control_s1_chipselect -> uart1_wr_control:chipselect
	wire         mm_interconnect_0_uart1_wr_control_s1_write;                 // mm_interconnect_0:uart1_wr_control_s1_write -> uart1_wr_control:write_n
	wire  [31:0] mm_interconnect_0_uart1_wr_control_s1_readdata;              // uart1_wr_control:readdata -> mm_interconnect_0:uart1_wr_control_s1_readdata
	wire         nios2e_instruction_master_waitrequest;                       // mm_interconnect_0:nios2e_instruction_master_waitrequest -> nios2e:i_waitrequest
	wire  [16:0] nios2e_instruction_master_address;                           // nios2e:i_address -> mm_interconnect_0:nios2e_instruction_master_address
	wire         nios2e_instruction_master_read;                              // nios2e:i_read -> mm_interconnect_0:nios2e_instruction_master_read
	wire  [31:0] nios2e_instruction_master_readdata;                          // mm_interconnect_0:nios2e_instruction_master_readdata -> nios2e:i_readdata
	wire  [31:0] mm_interconnect_0_onchip_ram_s1_writedata;                   // mm_interconnect_0:onchip_ram_s1_writedata -> onchip_ram:writedata
	wire  [13:0] mm_interconnect_0_onchip_ram_s1_address;                     // mm_interconnect_0:onchip_ram_s1_address -> onchip_ram:address
	wire         mm_interconnect_0_onchip_ram_s1_chipselect;                  // mm_interconnect_0:onchip_ram_s1_chipselect -> onchip_ram:chipselect
	wire         mm_interconnect_0_onchip_ram_s1_clken;                       // mm_interconnect_0:onchip_ram_s1_clken -> onchip_ram:clken
	wire         mm_interconnect_0_onchip_ram_s1_write;                       // mm_interconnect_0:onchip_ram_s1_write -> onchip_ram:write
	wire  [31:0] mm_interconnect_0_onchip_ram_s1_readdata;                    // onchip_ram:readdata -> mm_interconnect_0:onchip_ram_s1_readdata
	wire   [3:0] mm_interconnect_0_onchip_ram_s1_byteenable;                  // mm_interconnect_0:onchip_ram_s1_byteenable -> onchip_ram:byteenable
	wire         mm_interconnect_0_nios2e_jtag_debug_module_waitrequest;      // nios2e:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2e_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_nios2e_jtag_debug_module_writedata;        // mm_interconnect_0:nios2e_jtag_debug_module_writedata -> nios2e:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_nios2e_jtag_debug_module_address;          // mm_interconnect_0:nios2e_jtag_debug_module_address -> nios2e:jtag_debug_module_address
	wire         mm_interconnect_0_nios2e_jtag_debug_module_write;            // mm_interconnect_0:nios2e_jtag_debug_module_write -> nios2e:jtag_debug_module_write
	wire         mm_interconnect_0_nios2e_jtag_debug_module_read;             // mm_interconnect_0:nios2e_jtag_debug_module_read -> nios2e:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_nios2e_jtag_debug_module_readdata;         // nios2e:jtag_debug_module_readdata -> mm_interconnect_0:nios2e_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2e_jtag_debug_module_debugaccess;      // mm_interconnect_0:nios2e_jtag_debug_module_debugaccess -> nios2e:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_nios2e_jtag_debug_module_byteenable;       // mm_interconnect_0:nios2e_jtag_debug_module_byteenable -> nios2e:jtag_debug_module_byteenable
	wire   [1:0] mm_interconnect_0_sseg_counter_of_s1_address;                // mm_interconnect_0:sseg_counter_of_s1_address -> sseg_counter_of:address
	wire  [31:0] mm_interconnect_0_sseg_counter_of_s1_readdata;               // sseg_counter_of:readdata -> mm_interconnect_0:sseg_counter_of_s1_readdata
	wire   [1:0] mm_interconnect_0_leds1_counter_of_s1_address;               // mm_interconnect_0:leds1_counter_of_s1_address -> leds1_counter_of:address
	wire  [31:0] mm_interconnect_0_leds1_counter_of_s1_readdata;              // leds1_counter_of:readdata -> mm_interconnect_0:leds1_counter_of_s1_readdata
	wire  [31:0] mm_interconnect_0_bcd1_control_s1_writedata;                 // mm_interconnect_0:bcd1_control_s1_writedata -> bcd1_control:writedata
	wire   [1:0] mm_interconnect_0_bcd1_control_s1_address;                   // mm_interconnect_0:bcd1_control_s1_address -> bcd1_control:address
	wire         mm_interconnect_0_bcd1_control_s1_chipselect;                // mm_interconnect_0:bcd1_control_s1_chipselect -> bcd1_control:chipselect
	wire         mm_interconnect_0_bcd1_control_s1_write;                     // mm_interconnect_0:bcd1_control_s1_write -> bcd1_control:write_n
	wire  [31:0] mm_interconnect_0_bcd1_control_s1_readdata;                  // bcd1_control:readdata -> mm_interconnect_0:bcd1_control_s1_readdata
	wire  [31:0] mm_interconnect_0_rc1_ready_s1_writedata;                    // mm_interconnect_0:rc1_ready_s1_writedata -> rc1_ready:writedata
	wire   [1:0] mm_interconnect_0_rc1_ready_s1_address;                      // mm_interconnect_0:rc1_ready_s1_address -> rc1_ready:address
	wire         mm_interconnect_0_rc1_ready_s1_chipselect;                   // mm_interconnect_0:rc1_ready_s1_chipselect -> rc1_ready:chipselect
	wire         mm_interconnect_0_rc1_ready_s1_write;                        // mm_interconnect_0:rc1_ready_s1_write -> rc1_ready:write_n
	wire  [31:0] mm_interconnect_0_rc1_ready_s1_readdata;                     // rc1_ready:readdata -> mm_interconnect_0:rc1_ready_s1_readdata
	wire  [31:0] mm_interconnect_0_leds2_wr_val_s1_writedata;                 // mm_interconnect_0:leds2_wr_val_s1_writedata -> leds2_wr_val:writedata
	wire   [1:0] mm_interconnect_0_leds2_wr_val_s1_address;                   // mm_interconnect_0:leds2_wr_val_s1_address -> leds2_wr_val:address
	wire         mm_interconnect_0_leds2_wr_val_s1_chipselect;                // mm_interconnect_0:leds2_wr_val_s1_chipselect -> leds2_wr_val:chipselect
	wire         mm_interconnect_0_leds2_wr_val_s1_write;                     // mm_interconnect_0:leds2_wr_val_s1_write -> leds2_wr_val:write_n
	wire  [31:0] mm_interconnect_0_leds2_wr_val_s1_readdata;                  // leds2_wr_val:readdata -> mm_interconnect_0:leds2_wr_val_s1_readdata
	wire  [31:0] mm_interconnect_0_leds1_brightness_s1_writedata;             // mm_interconnect_0:leds1_brightness_s1_writedata -> leds1_brightness:writedata
	wire   [1:0] mm_interconnect_0_leds1_brightness_s1_address;               // mm_interconnect_0:leds1_brightness_s1_address -> leds1_brightness:address
	wire         mm_interconnect_0_leds1_brightness_s1_chipselect;            // mm_interconnect_0:leds1_brightness_s1_chipselect -> leds1_brightness:chipselect
	wire         mm_interconnect_0_leds1_brightness_s1_write;                 // mm_interconnect_0:leds1_brightness_s1_write -> leds1_brightness:write_n
	wire  [31:0] mm_interconnect_0_leds1_brightness_s1_readdata;              // leds1_brightness:readdata -> mm_interconnect_0:leds1_brightness_s1_readdata
	wire   [1:0] mm_interconnect_0_tc2_status_s1_address;                     // mm_interconnect_0:tc2_status_s1_address -> tc2_status:address
	wire  [31:0] mm_interconnect_0_tc2_status_s1_readdata;                    // tc2_status:readdata -> mm_interconnect_0:tc2_status_s1_readdata
	wire  [31:0] mm_interconnect_0_bcd1_bin_s1_writedata;                     // mm_interconnect_0:bcd1_bin_s1_writedata -> bcd1_bin:writedata
	wire   [1:0] mm_interconnect_0_bcd1_bin_s1_address;                       // mm_interconnect_0:bcd1_bin_s1_address -> bcd1_bin:address
	wire         mm_interconnect_0_bcd1_bin_s1_chipselect;                    // mm_interconnect_0:bcd1_bin_s1_chipselect -> bcd1_bin:chipselect
	wire         mm_interconnect_0_bcd1_bin_s1_write;                         // mm_interconnect_0:bcd1_bin_s1_write -> bcd1_bin:write_n
	wire  [31:0] mm_interconnect_0_bcd1_bin_s1_readdata;                      // bcd1_bin:readdata -> mm_interconnect_0:bcd1_bin_s1_readdata
	wire   [1:0] mm_interconnect_0_leds2_counter_of_s1_address;               // mm_interconnect_0:leds2_counter_of_s1_address -> leds2_counter_of:address
	wire  [31:0] mm_interconnect_0_leds2_counter_of_s1_readdata;              // leds2_counter_of:readdata -> mm_interconnect_0:leds2_counter_of_s1_readdata
	wire  [31:0] mm_interconnect_0_leds1_wr_val_s1_writedata;                 // mm_interconnect_0:leds1_wr_val_s1_writedata -> leds1_wr_val:writedata
	wire   [1:0] mm_interconnect_0_leds1_wr_val_s1_address;                   // mm_interconnect_0:leds1_wr_val_s1_address -> leds1_wr_val:address
	wire         mm_interconnect_0_leds1_wr_val_s1_chipselect;                // mm_interconnect_0:leds1_wr_val_s1_chipselect -> leds1_wr_val:chipselect
	wire         mm_interconnect_0_leds1_wr_val_s1_write;                     // mm_interconnect_0:leds1_wr_val_s1_write -> leds1_wr_val:write_n
	wire  [31:0] mm_interconnect_0_leds1_wr_val_s1_readdata;                  // leds1_wr_val:readdata -> mm_interconnect_0:leds1_wr_val_s1_readdata
	wire   [1:0] mm_interconnect_0_bcd1_bcd_s1_address;                       // mm_interconnect_0:bcd1_bcd_s1_address -> bcd1_bcd:address
	wire  [31:0] mm_interconnect_0_bcd1_bcd_s1_readdata;                      // bcd1_bcd:readdata -> mm_interconnect_0:bcd1_bcd_s1_readdata
	wire   [1:0] mm_interconnect_0_tc3_status_s1_address;                     // mm_interconnect_0:tc3_status_s1_address -> tc3_status:address
	wire  [31:0] mm_interconnect_0_tc3_status_s1_readdata;                    // tc3_status:readdata -> mm_interconnect_0:tc3_status_s1_readdata
	wire  [31:0] mm_interconnect_0_sseg_wr_val_s1_writedata;                  // mm_interconnect_0:sseg_wr_val_s1_writedata -> sseg_wr_val:writedata
	wire   [1:0] mm_interconnect_0_sseg_wr_val_s1_address;                    // mm_interconnect_0:sseg_wr_val_s1_address -> sseg_wr_val:address
	wire         mm_interconnect_0_sseg_wr_val_s1_chipselect;                 // mm_interconnect_0:sseg_wr_val_s1_chipselect -> sseg_wr_val:chipselect
	wire         mm_interconnect_0_sseg_wr_val_s1_write;                      // mm_interconnect_0:sseg_wr_val_s1_write -> sseg_wr_val:write_n
	wire  [31:0] mm_interconnect_0_sseg_wr_val_s1_readdata;                   // sseg_wr_val:readdata -> mm_interconnect_0:sseg_wr_val_s1_readdata
	wire  [31:0] mm_interconnect_0_sseg_brightness_s1_writedata;              // mm_interconnect_0:sseg_brightness_s1_writedata -> sseg_brightness:writedata
	wire   [1:0] mm_interconnect_0_sseg_brightness_s1_address;                // mm_interconnect_0:sseg_brightness_s1_address -> sseg_brightness:address
	wire         mm_interconnect_0_sseg_brightness_s1_chipselect;             // mm_interconnect_0:sseg_brightness_s1_chipselect -> sseg_brightness:chipselect
	wire         mm_interconnect_0_sseg_brightness_s1_write;                  // mm_interconnect_0:sseg_brightness_s1_write -> sseg_brightness:write_n
	wire  [31:0] mm_interconnect_0_sseg_brightness_s1_readdata;               // sseg_brightness:readdata -> mm_interconnect_0:sseg_brightness_s1_readdata
	wire  [31:0] mm_interconnect_0_uart1_dvsr_s1_writedata;                   // mm_interconnect_0:uart1_dvsr_s1_writedata -> uart1_dvsr:writedata
	wire   [1:0] mm_interconnect_0_uart1_dvsr_s1_address;                     // mm_interconnect_0:uart1_dvsr_s1_address -> uart1_dvsr:address
	wire         mm_interconnect_0_uart1_dvsr_s1_chipselect;                  // mm_interconnect_0:uart1_dvsr_s1_chipselect -> uart1_dvsr:chipselect
	wire         mm_interconnect_0_uart1_dvsr_s1_write;                       // mm_interconnect_0:uart1_dvsr_s1_write -> uart1_dvsr:write_n
	wire  [31:0] mm_interconnect_0_uart1_dvsr_s1_readdata;                    // uart1_dvsr:readdata -> mm_interconnect_0:uart1_dvsr_s1_readdata
	wire  [31:0] mm_interconnect_0_leds2_reset_control_s1_writedata;          // mm_interconnect_0:leds2_reset_control_s1_writedata -> leds2_reset_control:writedata
	wire   [1:0] mm_interconnect_0_leds2_reset_control_s1_address;            // mm_interconnect_0:leds2_reset_control_s1_address -> leds2_reset_control:address
	wire         mm_interconnect_0_leds2_reset_control_s1_chipselect;         // mm_interconnect_0:leds2_reset_control_s1_chipselect -> leds2_reset_control:chipselect
	wire         mm_interconnect_0_leds2_reset_control_s1_write;              // mm_interconnect_0:leds2_reset_control_s1_write -> leds2_reset_control:write_n
	wire  [31:0] mm_interconnect_0_leds2_reset_control_s1_readdata;           // leds2_reset_control:readdata -> mm_interconnect_0:leds2_reset_control_s1_readdata
	wire  [31:0] mm_interconnect_0_warn_pwm_brightness_s1_writedata;          // mm_interconnect_0:warn_pwm_brightness_s1_writedata -> warn_pwm_brightness:writedata
	wire   [1:0] mm_interconnect_0_warn_pwm_brightness_s1_address;            // mm_interconnect_0:warn_pwm_brightness_s1_address -> warn_pwm_brightness:address
	wire         mm_interconnect_0_warn_pwm_brightness_s1_chipselect;         // mm_interconnect_0:warn_pwm_brightness_s1_chipselect -> warn_pwm_brightness:chipselect
	wire         mm_interconnect_0_warn_pwm_brightness_s1_write;              // mm_interconnect_0:warn_pwm_brightness_s1_write -> warn_pwm_brightness:write_n
	wire  [31:0] mm_interconnect_0_warn_pwm_brightness_s1_readdata;           // warn_pwm_brightness:readdata -> mm_interconnect_0:warn_pwm_brightness_s1_readdata
	wire   [1:0] mm_interconnect_0_bcd1_status_s1_address;                    // mm_interconnect_0:bcd1_status_s1_address -> bcd1_status:address
	wire  [31:0] mm_interconnect_0_bcd1_status_s1_readdata;                   // bcd1_status:readdata -> mm_interconnect_0:bcd1_status_s1_readdata
	wire  [31:0] mm_interconnect_0_daylight_s1_writedata;                     // mm_interconnect_0:daylight_s1_writedata -> daylight:writedata
	wire   [1:0] mm_interconnect_0_daylight_s1_address;                       // mm_interconnect_0:daylight_s1_address -> daylight:address
	wire         mm_interconnect_0_daylight_s1_chipselect;                    // mm_interconnect_0:daylight_s1_chipselect -> daylight:chipselect
	wire         mm_interconnect_0_daylight_s1_write;                         // mm_interconnect_0:daylight_s1_write -> daylight:write_n
	wire  [31:0] mm_interconnect_0_daylight_s1_readdata;                      // daylight:readdata -> mm_interconnect_0:daylight_s1_readdata
	wire  [31:0] mm_interconnect_0_uart1_baud_control_s1_writedata;           // mm_interconnect_0:uart1_baud_control_s1_writedata -> uart1_baud_control:writedata
	wire   [1:0] mm_interconnect_0_uart1_baud_control_s1_address;             // mm_interconnect_0:uart1_baud_control_s1_address -> uart1_baud_control:address
	wire         mm_interconnect_0_uart1_baud_control_s1_chipselect;          // mm_interconnect_0:uart1_baud_control_s1_chipselect -> uart1_baud_control:chipselect
	wire         mm_interconnect_0_uart1_baud_control_s1_write;               // mm_interconnect_0:uart1_baud_control_s1_write -> uart1_baud_control:write_n
	wire  [31:0] mm_interconnect_0_uart1_baud_control_s1_readdata;            // uart1_baud_control:readdata -> mm_interconnect_0:uart1_baud_control_s1_readdata
	wire   [1:0] mm_interconnect_0_bcd1_counter_s1_address;                   // mm_interconnect_0:bcd1_counter_s1_address -> bcd1_counter:address
	wire  [31:0] mm_interconnect_0_bcd1_counter_s1_readdata;                  // bcd1_counter:readdata -> mm_interconnect_0:bcd1_counter_s1_readdata
	wire  [31:0] mm_interconnect_0_led_period_s1_writedata;                   // mm_interconnect_0:led_period_s1_writedata -> led_period:writedata
	wire   [1:0] mm_interconnect_0_led_period_s1_address;                     // mm_interconnect_0:led_period_s1_address -> led_period:address
	wire         mm_interconnect_0_led_period_s1_chipselect;                  // mm_interconnect_0:led_period_s1_chipselect -> led_period:chipselect
	wire         mm_interconnect_0_led_period_s1_write;                       // mm_interconnect_0:led_period_s1_write -> led_period:write_n
	wire  [31:0] mm_interconnect_0_led_period_s1_readdata;                    // led_period:readdata -> mm_interconnect_0:led_period_s1_readdata
	wire   [0:0] mm_interconnect_0_sysid_c001_control_slave_address;          // mm_interconnect_0:sysid_c001_control_slave_address -> sysid_c001:address
	wire  [31:0] mm_interconnect_0_sysid_c001_control_slave_readdata;         // sysid_c001:readdata -> mm_interconnect_0:sysid_c001_control_slave_readdata
	wire  [31:0] mm_interconnect_0_status_led_en_s1_writedata;                // mm_interconnect_0:status_led_en_s1_writedata -> status_led_en:writedata
	wire   [2:0] mm_interconnect_0_status_led_en_s1_address;                  // mm_interconnect_0:status_led_en_s1_address -> status_led_en:address
	wire         mm_interconnect_0_status_led_en_s1_chipselect;               // mm_interconnect_0:status_led_en_s1_chipselect -> status_led_en:chipselect
	wire         mm_interconnect_0_status_led_en_s1_write;                    // mm_interconnect_0:status_led_en_s1_write -> status_led_en:write_n
	wire  [31:0] mm_interconnect_0_status_led_en_s1_readdata;                 // status_led_en:readdata -> mm_interconnect_0:status_led_en_s1_readdata
	wire  [31:0] mm_interconnect_0_tc2_m_s1_writedata;                        // mm_interconnect_0:tc2_m_s1_writedata -> tc2_m:writedata
	wire   [1:0] mm_interconnect_0_tc2_m_s1_address;                          // mm_interconnect_0:tc2_m_s1_address -> tc2_m:address
	wire         mm_interconnect_0_tc2_m_s1_chipselect;                       // mm_interconnect_0:tc2_m_s1_chipselect -> tc2_m:chipselect
	wire         mm_interconnect_0_tc2_m_s1_write;                            // mm_interconnect_0:tc2_m_s1_write -> tc2_m:write_n
	wire  [31:0] mm_interconnect_0_tc2_m_s1_readdata;                         // tc2_m:readdata -> mm_interconnect_0:tc2_m_s1_readdata
	wire   [1:0] mm_interconnect_0_uart1_tx_counter_s1_address;               // mm_interconnect_0:uart1_tx_counter_s1_address -> uart1_tx_counter:address
	wire  [31:0] mm_interconnect_0_uart1_tx_counter_s1_readdata;              // uart1_tx_counter:readdata -> mm_interconnect_0:uart1_tx_counter_s1_readdata
	wire   [1:0] mm_interconnect_0_uart1_r_data_s1_address;                   // mm_interconnect_0:uart1_r_data_s1_address -> uart1_r_data:address
	wire  [31:0] mm_interconnect_0_uart1_r_data_s1_readdata;                  // uart1_r_data:readdata -> mm_interconnect_0:uart1_r_data_s1_readdata
	wire  [31:0] mm_interconnect_0_tc1_m_s1_writedata;                        // mm_interconnect_0:tc1_m_s1_writedata -> tc1_m:writedata
	wire   [1:0] mm_interconnect_0_tc1_m_s1_address;                          // mm_interconnect_0:tc1_m_s1_address -> tc1_m:address
	wire         mm_interconnect_0_tc1_m_s1_chipselect;                       // mm_interconnect_0:tc1_m_s1_chipselect -> tc1_m:chipselect
	wire         mm_interconnect_0_tc1_m_s1_write;                            // mm_interconnect_0:tc1_m_s1_write -> tc1_m:write_n
	wire  [31:0] mm_interconnect_0_tc1_m_s1_readdata;                         // tc1_m:readdata -> mm_interconnect_0:tc1_m_s1_readdata
	wire         nios2e_data_master_waitrequest;                              // mm_interconnect_0:nios2e_data_master_waitrequest -> nios2e:d_waitrequest
	wire  [31:0] nios2e_data_master_writedata;                                // nios2e:d_writedata -> mm_interconnect_0:nios2e_data_master_writedata
	wire  [16:0] nios2e_data_master_address;                                  // nios2e:d_address -> mm_interconnect_0:nios2e_data_master_address
	wire         nios2e_data_master_write;                                    // nios2e:d_write -> mm_interconnect_0:nios2e_data_master_write
	wire         nios2e_data_master_read;                                     // nios2e:d_read -> mm_interconnect_0:nios2e_data_master_read
	wire  [31:0] nios2e_data_master_readdata;                                 // mm_interconnect_0:nios2e_data_master_readdata -> nios2e:d_readdata
	wire         nios2e_data_master_debugaccess;                              // nios2e:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2e_data_master_debugaccess
	wire   [3:0] nios2e_data_master_byteenable;                               // nios2e:d_byteenable -> mm_interconnect_0:nios2e_data_master_byteenable
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire  [31:0] mm_interconnect_0_leds2_brightness_s1_writedata;             // mm_interconnect_0:leds2_brightness_s1_writedata -> leds2_brightness:writedata
	wire   [1:0] mm_interconnect_0_leds2_brightness_s1_address;               // mm_interconnect_0:leds2_brightness_s1_address -> leds2_brightness:address
	wire         mm_interconnect_0_leds2_brightness_s1_chipselect;            // mm_interconnect_0:leds2_brightness_s1_chipselect -> leds2_brightness:chipselect
	wire         mm_interconnect_0_leds2_brightness_s1_write;                 // mm_interconnect_0:leds2_brightness_s1_write -> leds2_brightness:write_n
	wire  [31:0] mm_interconnect_0_leds2_brightness_s1_readdata;              // leds2_brightness:readdata -> mm_interconnect_0:leds2_brightness_s1_readdata
	wire   [1:0] mm_interconnect_0_sseg_counter_s1_address;                   // mm_interconnect_0:sseg_counter_s1_address -> sseg_counter:address
	wire  [31:0] mm_interconnect_0_sseg_counter_s1_readdata;                  // sseg_counter:readdata -> mm_interconnect_0:sseg_counter_s1_readdata
	wire  [31:0] mm_interconnect_0_uart1_reset_control_s1_writedata;          // mm_interconnect_0:uart1_reset_control_s1_writedata -> uart1_reset_control:writedata
	wire   [1:0] mm_interconnect_0_uart1_reset_control_s1_address;            // mm_interconnect_0:uart1_reset_control_s1_address -> uart1_reset_control:address
	wire         mm_interconnect_0_uart1_reset_control_s1_chipselect;         // mm_interconnect_0:uart1_reset_control_s1_chipselect -> uart1_reset_control:chipselect
	wire         mm_interconnect_0_uart1_reset_control_s1_write;              // mm_interconnect_0:uart1_reset_control_s1_write -> uart1_reset_control:write_n
	wire  [31:0] mm_interconnect_0_uart1_reset_control_s1_readdata;           // uart1_reset_control:readdata -> mm_interconnect_0:uart1_reset_control_s1_readdata
	wire  [31:0] mm_interconnect_0_sseg_reset_control_s1_writedata;           // mm_interconnect_0:sseg_reset_control_s1_writedata -> sseg_reset_control:writedata
	wire   [1:0] mm_interconnect_0_sseg_reset_control_s1_address;             // mm_interconnect_0:sseg_reset_control_s1_address -> sseg_reset_control:address
	wire         mm_interconnect_0_sseg_reset_control_s1_chipselect;          // mm_interconnect_0:sseg_reset_control_s1_chipselect -> sseg_reset_control:chipselect
	wire         mm_interconnect_0_sseg_reset_control_s1_write;               // mm_interconnect_0:sseg_reset_control_s1_write -> sseg_reset_control:write_n
	wire  [31:0] mm_interconnect_0_sseg_reset_control_s1_readdata;            // sseg_reset_control:readdata -> mm_interconnect_0:sseg_reset_control_s1_readdata
	wire  [31:0] mm_interconnect_0_warn_pwm_control_s1_writedata;             // mm_interconnect_0:warn_pwm_control_s1_writedata -> warn_pwm_control:writedata
	wire   [1:0] mm_interconnect_0_warn_pwm_control_s1_address;               // mm_interconnect_0:warn_pwm_control_s1_address -> warn_pwm_control:address
	wire         mm_interconnect_0_warn_pwm_control_s1_chipselect;            // mm_interconnect_0:warn_pwm_control_s1_chipselect -> warn_pwm_control:chipselect
	wire         mm_interconnect_0_warn_pwm_control_s1_write;                 // mm_interconnect_0:warn_pwm_control_s1_write -> warn_pwm_control:write_n
	wire  [31:0] mm_interconnect_0_warn_pwm_control_s1_readdata;              // warn_pwm_control:readdata -> mm_interconnect_0:warn_pwm_control_s1_readdata
	wire   [1:0] mm_interconnect_0_leds1_counter_s1_address;                  // mm_interconnect_0:leds1_counter_s1_address -> leds1_counter:address
	wire  [31:0] mm_interconnect_0_leds1_counter_s1_readdata;                 // leds1_counter:readdata -> mm_interconnect_0:leds1_counter_s1_readdata
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // rc1_ready:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                    // daylight:irq -> irq_mapper:receiver2_irq
	wire  [31:0] nios2e_d_irq_irq;                                            // irq_mapper:sender_irq -> nios2e:d_irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [bcd1_bcd:reset_n, bcd1_bin:reset_n, bcd1_control:reset_n, bcd1_counter:reset_n, bcd1_status:reset_n, daylight:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, led_period:reset_n, leds1_brightness:reset_n, leds1_counter:reset_n, leds1_counter_of:reset_n, leds1_reset_control:reset_n, leds1_wr_val:reset_n, leds2_brightness:reset_n, leds2_counter:reset_n, leds2_counter_of:reset_n, leds2_reset_control:reset_n, leds2_wr_val:reset_n, mm_interconnect_0:nios2e_reset_n_reset_bridge_in_reset_reset, nios2e:reset_n, onchip_ram:reset, rc1_control:reset_n, rc1_ready:reset_n, rst_translator:in_reset, sseg_brightness:reset_n, sseg_counter:reset_n, sseg_counter_of:reset_n, sseg_reset_control:reset_n, sseg_wr_val:reset_n, status_led_en:reset_n, sysid_c001:reset_n, tc1_m:reset_n, tc1_status:reset_n, tc2_m:reset_n, tc2_status:reset_n, tc3_m:reset_n, tc3_status:reset_n, tc4_m:reset_n, tc4_status:reset_n, tc_reset_control:reset_n, uart1_baud_control:reset_n, uart1_dvsr:reset_n, uart1_r_data:reset_n, uart1_reset_control:reset_n, uart1_rx_counter:reset_n, uart1_status_control:reset_n, uart1_tx_counter:reset_n, uart1_w_data:reset_n, uart1_wr_control:reset_n, warn_pwm_brightness:reset_n, warn_pwm_control:reset_n]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [nios2e:reset_req, onchip_ram:reset_req, rst_translator:reset_req_in]
	wire         nios2e_jtag_debug_module_reset_reset;                        // nios2e:jtag_debug_module_resetrequest -> rst_controller:reset_in1

	controller_sysid_c001 sysid_c001 (
		.clock    (clock_50_clk),                                        //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                     //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_c001_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_c001_control_slave_address)   //              .address
	);

	controller_jtag_uart_0 jtag_uart_0 (
		.clk            (clock_50_clk),                                                //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	controller_nios2e nios2e (
		.clk                                   (clock_50_clk),                                           //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                        //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                     //                          .reset_req
		.d_address                             (nios2e_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2e_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2e_data_master_read),                                //                          .read
		.d_readdata                            (nios2e_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2e_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2e_data_master_write),                               //                          .write
		.d_writedata                           (nios2e_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios2e_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2e_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2e_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2e_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2e_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (nios2e_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2e_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2e_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2e_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2e_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2e_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2e_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2e_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2e_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2e_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                        // custom_instruction_master.readra
	);

	controller_onchip_ram onchip_ram (
		.clk        (clock_50_clk),                               //   clk1.clk
		.address    (mm_interconnect_0_onchip_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)          //       .reset_req
	);

	controller_daylight daylight (
		.clk        (clock_50_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_daylight_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_daylight_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_daylight_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_daylight_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_daylight_s1_readdata),   //                    .readdata
		.in_port    (daylight_export),                          // external_connection.export
		.irq        (irq_mapper_receiver2_irq)                  //                 irq.irq
	);

	controller_tc1_m tc1_m (
		.clk        (clock_50_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_tc1_m_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_tc1_m_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_tc1_m_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_tc1_m_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_tc1_m_s1_readdata),   //                    .readdata
		.out_port   (tc1_m_export)                           // external_connection.export
	);

	controller_tc1_m tc2_m (
		.clk        (clock_50_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_tc2_m_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_tc2_m_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_tc2_m_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_tc2_m_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_tc2_m_s1_readdata),   //                    .readdata
		.out_port   (tc2_m_export)                           // external_connection.export
	);

	controller_tc1_m tc3_m (
		.clk        (clock_50_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_tc3_m_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_tc3_m_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_tc3_m_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_tc3_m_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_tc3_m_s1_readdata),   //                    .readdata
		.out_port   (tc3_m_export)                           // external_connection.export
	);

	controller_tc1_m tc4_m (
		.clk        (clock_50_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_tc4_m_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_tc4_m_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_tc4_m_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_tc4_m_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_tc4_m_s1_readdata),   //                    .readdata
		.out_port   (tc4_m_export)                           // external_connection.export
	);

	controller_tc_reset_control tc_reset_control (
		.clk        (clock_50_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_0_tc_reset_control_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_tc_reset_control_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_tc_reset_control_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_tc_reset_control_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_tc_reset_control_s1_readdata),   //                    .readdata
		.out_port   (tc_reset_control_export)                           // external_connection.export
	);

	controller_tc1_status tc1_status (
		.clk      (clock_50_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_tc1_status_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_tc1_status_s1_readdata), //                    .readdata
		.in_port  (tc1_status_export)                         // external_connection.export
	);

	controller_tc1_status tc2_status (
		.clk      (clock_50_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_tc2_status_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_tc2_status_s1_readdata), //                    .readdata
		.in_port  (tc2_status_export)                         // external_connection.export
	);

	controller_tc1_status tc3_status (
		.clk      (clock_50_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_tc3_status_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_tc3_status_s1_readdata), //                    .readdata
		.in_port  (tc3_status_export)                         // external_connection.export
	);

	controller_tc1_status tc4_status (
		.clk      (clock_50_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_tc4_status_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_tc4_status_s1_readdata), //                    .readdata
		.in_port  (tc4_status_export)                         // external_connection.export
	);

	controller_uart1_w_data uart1_w_data (
		.clk        (clock_50_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_uart1_w_data_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_uart1_w_data_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_uart1_w_data_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_uart1_w_data_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_uart1_w_data_s1_readdata),   //                    .readdata
		.out_port   (uart1_w_data_export)                           // external_connection.export
	);

	controller_uart1_reset_control uart1_reset_control (
		.clk        (clock_50_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                     //               reset.reset_n
		.address    (mm_interconnect_0_uart1_reset_control_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_uart1_reset_control_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_uart1_reset_control_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_uart1_reset_control_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_uart1_reset_control_s1_readdata),   //                    .readdata
		.out_port   (uart1_reset_control_export)                           // external_connection.export
	);

	controller_uart1_wr_control uart1_wr_control (
		.clk        (clock_50_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_0_uart1_wr_control_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_uart1_wr_control_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_uart1_wr_control_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_uart1_wr_control_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_uart1_wr_control_s1_readdata),   //                    .readdata
		.out_port   (uart1_wr_control_export)                           // external_connection.export
	);

	controller_uart1_baud_control uart1_baud_control (
		.clk        (clock_50_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                    //               reset.reset_n
		.address    (mm_interconnect_0_uart1_baud_control_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_uart1_baud_control_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_uart1_baud_control_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_uart1_baud_control_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_uart1_baud_control_s1_readdata),   //                    .readdata
		.out_port   (uart1_baud_control_export)                           // external_connection.export
	);

	controller_uart1_r_data uart1_r_data (
		.clk      (clock_50_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_0_uart1_r_data_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_uart1_r_data_s1_readdata), //                    .readdata
		.in_port  (uart1_r_data_export)                         // external_connection.export
	);

	controller_uart1_r_data uart1_rx_counter (
		.clk      (clock_50_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address  (mm_interconnect_0_uart1_rx_counter_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_uart1_rx_counter_s1_readdata), //                    .readdata
		.in_port  (uart1_rx_counter_export)                         // external_connection.export
	);

	controller_uart1_r_data uart1_tx_counter (
		.clk      (clock_50_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address  (mm_interconnect_0_uart1_tx_counter_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_uart1_tx_counter_s1_readdata), //                    .readdata
		.in_port  (uart1_tx_counter_export)                         // external_connection.export
	);

	controller_uart1_status_control uart1_status_control (
		.clk      (clock_50_clk),                                       //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                    //               reset.reset_n
		.address  (mm_interconnect_0_uart1_status_control_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_uart1_status_control_s1_readdata), //                    .readdata
		.in_port  (uart1_status_control_export)                         // external_connection.export
	);

	controller_bcd1_bin bcd1_bin (
		.clk        (clock_50_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_bcd1_bin_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bcd1_bin_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bcd1_bin_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bcd1_bin_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bcd1_bin_s1_readdata),   //                    .readdata
		.out_port   (bcd1_bin_export)                           // external_connection.export
	);

	controller_bcd1_control bcd1_control (
		.clk        (clock_50_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_bcd1_control_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bcd1_control_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bcd1_control_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bcd1_control_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bcd1_control_s1_readdata),   //                    .readdata
		.out_port   (bcd1_control_export)                           // external_connection.export
	);

	controller_bcd1_bcd bcd1_bcd (
		.clk      (clock_50_clk),                           //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_bcd1_bcd_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_bcd1_bcd_s1_readdata), //                    .readdata
		.in_port  (bcd1_bcd_export)                         // external_connection.export
	);

	controller_uart1_r_data bcd1_counter (
		.clk      (clock_50_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_0_bcd1_counter_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_bcd1_counter_s1_readdata), //                    .readdata
		.in_port  (bcd1_counter_export)                         // external_connection.export
	);

	controller_bcd1_status bcd1_status (
		.clk      (clock_50_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_bcd1_status_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_bcd1_status_s1_readdata), //                    .readdata
		.in_port  (bcd1_status_export)                         // external_connection.export
	);

	controller_uart1_w_data warn_pwm_brightness (
		.clk        (clock_50_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                     //               reset.reset_n
		.address    (mm_interconnect_0_warn_pwm_brightness_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_warn_pwm_brightness_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_warn_pwm_brightness_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_warn_pwm_brightness_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_warn_pwm_brightness_s1_readdata),   //                    .readdata
		.out_port   (warn_pwm_brightness_export)                           // external_connection.export
	);

	controller_status_led_en status_led_en (
		.clk        (clock_50_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_status_led_en_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_status_led_en_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_status_led_en_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_status_led_en_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_status_led_en_s1_readdata),   //                    .readdata
		.out_port   (status_led_en_export)                           // external_connection.export
	);

	controller_warn_pwm_control warn_pwm_control (
		.clk        (clock_50_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_0_warn_pwm_control_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_warn_pwm_control_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_warn_pwm_control_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_warn_pwm_control_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_warn_pwm_control_s1_readdata),   //                    .readdata
		.out_port   (warn_pwm_control_export)                           // external_connection.export
	);

	controller_uart1_w_data sseg_brightness (
		.clk        (clock_50_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_sseg_brightness_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sseg_brightness_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sseg_brightness_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sseg_brightness_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sseg_brightness_s1_readdata),   //                    .readdata
		.out_port   (sseg_brightness_export)                           // external_connection.export
	);

	controller_sseg_reset_control sseg_reset_control (
		.clk        (clock_50_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                    //               reset.reset_n
		.address    (mm_interconnect_0_sseg_reset_control_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sseg_reset_control_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sseg_reset_control_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sseg_reset_control_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sseg_reset_control_s1_readdata),   //                    .readdata
		.out_port   (sseg_reset_control_export)                           // external_connection.export
	);

	controller_sseg_wr_val sseg_wr_val (
		.clk        (clock_50_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_sseg_wr_val_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sseg_wr_val_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sseg_wr_val_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sseg_wr_val_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sseg_wr_val_s1_readdata),   //                    .readdata
		.out_port   (sseg_wr_val_export)                           // external_connection.export
	);

	controller_uart1_r_data sseg_counter (
		.clk      (clock_50_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_0_sseg_counter_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_sseg_counter_s1_readdata), //                    .readdata
		.in_port  (sseg_counter_export)                         // external_connection.export
	);

	controller_sseg_counter_of sseg_counter_of (
		.clk      (clock_50_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address  (mm_interconnect_0_sseg_counter_of_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_sseg_counter_of_s1_readdata), //                    .readdata
		.in_port  (sseg_counter_of_export)                         // external_connection.export
	);

	controller_uart1_w_data leds1_brightness (
		.clk        (clock_50_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_0_leds1_brightness_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds1_brightness_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds1_brightness_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds1_brightness_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds1_brightness_s1_readdata),   //                    .readdata
		.out_port   (leds1_brightness_export)                           // external_connection.export
	);

	controller_sseg_reset_control leds1_reset_control (
		.clk        (clock_50_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                     //               reset.reset_n
		.address    (mm_interconnect_0_leds1_reset_control_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds1_reset_control_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds1_reset_control_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds1_reset_control_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds1_reset_control_s1_readdata),   //                    .readdata
		.out_port   (leds1_reset_control_export)                           // external_connection.export
	);

	controller_leds1_wr_val leds1_wr_val (
		.clk        (clock_50_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_leds1_wr_val_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds1_wr_val_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds1_wr_val_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds1_wr_val_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds1_wr_val_s1_readdata),   //                    .readdata
		.out_port   (leds1_wr_val_export)                           // external_connection.export
	);

	controller_uart1_r_data leds1_counter (
		.clk      (clock_50_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address  (mm_interconnect_0_leds1_counter_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_leds1_counter_s1_readdata), //                    .readdata
		.in_port  (leds1_counter_export)                         // external_connection.export
	);

	controller_sseg_counter_of leds1_counter_of (
		.clk      (clock_50_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address  (mm_interconnect_0_leds1_counter_of_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_leds1_counter_of_s1_readdata), //                    .readdata
		.in_port  (leds1_counter_of_export)                         // external_connection.export
	);

	controller_uart1_dvsr uart1_dvsr (
		.clk        (clock_50_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_uart1_dvsr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_uart1_dvsr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_uart1_dvsr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_uart1_dvsr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_uart1_dvsr_s1_readdata),   //                    .readdata
		.out_port   (uart1_dvsr_export)                           // external_connection.export
	);

	controller_rc1_control rc1_control (
		.clk        (clock_50_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_rc1_control_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_rc1_control_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_rc1_control_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_rc1_control_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_rc1_control_s1_readdata),   //                    .readdata
		.out_port   (rc1_control_export)                           // external_connection.export
	);

	controller_daylight rc1_ready (
		.clk        (clock_50_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_rc1_ready_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_rc1_ready_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_rc1_ready_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_rc1_ready_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_rc1_ready_s1_readdata),   //                    .readdata
		.in_port    (rc1_ready_export),                          // external_connection.export
		.irq        (irq_mapper_receiver1_irq)                   //                 irq.irq
	);

	controller_led_period led_period (
		.clk        (clock_50_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_led_period_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_period_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_period_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_period_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_period_s1_readdata),   //                    .readdata
		.out_port   (led_period_export)                           // external_connection.export
	);

	controller_sseg_reset_control leds2_reset_control (
		.clk        (clock_50_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                     //               reset.reset_n
		.address    (mm_interconnect_0_leds2_reset_control_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds2_reset_control_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds2_reset_control_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds2_reset_control_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds2_reset_control_s1_readdata),   //                    .readdata
		.out_port   (leds2_reset_control_export)                           // external_connection.export
	);

	controller_leds1_wr_val leds2_wr_val (
		.clk        (clock_50_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_leds2_wr_val_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds2_wr_val_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds2_wr_val_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds2_wr_val_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds2_wr_val_s1_readdata),   //                    .readdata
		.out_port   (leds2_wr_val_export)                           // external_connection.export
	);

	controller_uart1_r_data leds2_counter (
		.clk      (clock_50_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address  (mm_interconnect_0_leds2_counter_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_leds2_counter_s1_readdata), //                    .readdata
		.in_port  (leds2_counter_export)                         // external_connection.export
	);

	controller_sseg_counter_of leds2_counter_of (
		.clk      (clock_50_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address  (mm_interconnect_0_leds2_counter_of_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_leds2_counter_of_s1_readdata), //                    .readdata
		.in_port  (leds2_counter_of_export)                         // external_connection.export
	);

	controller_uart1_w_data leds2_brightness (
		.clk        (clock_50_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_0_leds2_brightness_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds2_brightness_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds2_brightness_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds2_brightness_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds2_brightness_s1_readdata),   //                    .readdata
		.out_port   (leds2_brightness_export)                           // external_connection.export
	);

	controller_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                              (clock_50_clk),                                                //                            clk_0_clk.clk
		.nios2e_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                              // nios2e_reset_n_reset_bridge_in_reset.reset
		.nios2e_data_master_address                 (nios2e_data_master_address),                                  //                   nios2e_data_master.address
		.nios2e_data_master_waitrequest             (nios2e_data_master_waitrequest),                              //                                     .waitrequest
		.nios2e_data_master_byteenable              (nios2e_data_master_byteenable),                               //                                     .byteenable
		.nios2e_data_master_read                    (nios2e_data_master_read),                                     //                                     .read
		.nios2e_data_master_readdata                (nios2e_data_master_readdata),                                 //                                     .readdata
		.nios2e_data_master_write                   (nios2e_data_master_write),                                    //                                     .write
		.nios2e_data_master_writedata               (nios2e_data_master_writedata),                                //                                     .writedata
		.nios2e_data_master_debugaccess             (nios2e_data_master_debugaccess),                              //                                     .debugaccess
		.nios2e_instruction_master_address          (nios2e_instruction_master_address),                           //            nios2e_instruction_master.address
		.nios2e_instruction_master_waitrequest      (nios2e_instruction_master_waitrequest),                       //                                     .waitrequest
		.nios2e_instruction_master_read             (nios2e_instruction_master_read),                              //                                     .read
		.nios2e_instruction_master_readdata         (nios2e_instruction_master_readdata),                          //                                     .readdata
		.bcd1_bcd_s1_address                        (mm_interconnect_0_bcd1_bcd_s1_address),                       //                          bcd1_bcd_s1.address
		.bcd1_bcd_s1_readdata                       (mm_interconnect_0_bcd1_bcd_s1_readdata),                      //                                     .readdata
		.bcd1_bin_s1_address                        (mm_interconnect_0_bcd1_bin_s1_address),                       //                          bcd1_bin_s1.address
		.bcd1_bin_s1_write                          (mm_interconnect_0_bcd1_bin_s1_write),                         //                                     .write
		.bcd1_bin_s1_readdata                       (mm_interconnect_0_bcd1_bin_s1_readdata),                      //                                     .readdata
		.bcd1_bin_s1_writedata                      (mm_interconnect_0_bcd1_bin_s1_writedata),                     //                                     .writedata
		.bcd1_bin_s1_chipselect                     (mm_interconnect_0_bcd1_bin_s1_chipselect),                    //                                     .chipselect
		.bcd1_control_s1_address                    (mm_interconnect_0_bcd1_control_s1_address),                   //                      bcd1_control_s1.address
		.bcd1_control_s1_write                      (mm_interconnect_0_bcd1_control_s1_write),                     //                                     .write
		.bcd1_control_s1_readdata                   (mm_interconnect_0_bcd1_control_s1_readdata),                  //                                     .readdata
		.bcd1_control_s1_writedata                  (mm_interconnect_0_bcd1_control_s1_writedata),                 //                                     .writedata
		.bcd1_control_s1_chipselect                 (mm_interconnect_0_bcd1_control_s1_chipselect),                //                                     .chipselect
		.bcd1_counter_s1_address                    (mm_interconnect_0_bcd1_counter_s1_address),                   //                      bcd1_counter_s1.address
		.bcd1_counter_s1_readdata                   (mm_interconnect_0_bcd1_counter_s1_readdata),                  //                                     .readdata
		.bcd1_status_s1_address                     (mm_interconnect_0_bcd1_status_s1_address),                    //                       bcd1_status_s1.address
		.bcd1_status_s1_readdata                    (mm_interconnect_0_bcd1_status_s1_readdata),                   //                                     .readdata
		.daylight_s1_address                        (mm_interconnect_0_daylight_s1_address),                       //                          daylight_s1.address
		.daylight_s1_write                          (mm_interconnect_0_daylight_s1_write),                         //                                     .write
		.daylight_s1_readdata                       (mm_interconnect_0_daylight_s1_readdata),                      //                                     .readdata
		.daylight_s1_writedata                      (mm_interconnect_0_daylight_s1_writedata),                     //                                     .writedata
		.daylight_s1_chipselect                     (mm_interconnect_0_daylight_s1_chipselect),                    //                                     .chipselect
		.jtag_uart_0_avalon_jtag_slave_address      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //        jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                     .write
		.jtag_uart_0_avalon_jtag_slave_read         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                     .read
		.jtag_uart_0_avalon_jtag_slave_readdata     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                     .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                     .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                     .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                     .chipselect
		.led_period_s1_address                      (mm_interconnect_0_led_period_s1_address),                     //                        led_period_s1.address
		.led_period_s1_write                        (mm_interconnect_0_led_period_s1_write),                       //                                     .write
		.led_period_s1_readdata                     (mm_interconnect_0_led_period_s1_readdata),                    //                                     .readdata
		.led_period_s1_writedata                    (mm_interconnect_0_led_period_s1_writedata),                   //                                     .writedata
		.led_period_s1_chipselect                   (mm_interconnect_0_led_period_s1_chipselect),                  //                                     .chipselect
		.leds1_brightness_s1_address                (mm_interconnect_0_leds1_brightness_s1_address),               //                  leds1_brightness_s1.address
		.leds1_brightness_s1_write                  (mm_interconnect_0_leds1_brightness_s1_write),                 //                                     .write
		.leds1_brightness_s1_readdata               (mm_interconnect_0_leds1_brightness_s1_readdata),              //                                     .readdata
		.leds1_brightness_s1_writedata              (mm_interconnect_0_leds1_brightness_s1_writedata),             //                                     .writedata
		.leds1_brightness_s1_chipselect             (mm_interconnect_0_leds1_brightness_s1_chipselect),            //                                     .chipselect
		.leds1_counter_s1_address                   (mm_interconnect_0_leds1_counter_s1_address),                  //                     leds1_counter_s1.address
		.leds1_counter_s1_readdata                  (mm_interconnect_0_leds1_counter_s1_readdata),                 //                                     .readdata
		.leds1_counter_of_s1_address                (mm_interconnect_0_leds1_counter_of_s1_address),               //                  leds1_counter_of_s1.address
		.leds1_counter_of_s1_readdata               (mm_interconnect_0_leds1_counter_of_s1_readdata),              //                                     .readdata
		.leds1_reset_control_s1_address             (mm_interconnect_0_leds1_reset_control_s1_address),            //               leds1_reset_control_s1.address
		.leds1_reset_control_s1_write               (mm_interconnect_0_leds1_reset_control_s1_write),              //                                     .write
		.leds1_reset_control_s1_readdata            (mm_interconnect_0_leds1_reset_control_s1_readdata),           //                                     .readdata
		.leds1_reset_control_s1_writedata           (mm_interconnect_0_leds1_reset_control_s1_writedata),          //                                     .writedata
		.leds1_reset_control_s1_chipselect          (mm_interconnect_0_leds1_reset_control_s1_chipselect),         //                                     .chipselect
		.leds1_wr_val_s1_address                    (mm_interconnect_0_leds1_wr_val_s1_address),                   //                      leds1_wr_val_s1.address
		.leds1_wr_val_s1_write                      (mm_interconnect_0_leds1_wr_val_s1_write),                     //                                     .write
		.leds1_wr_val_s1_readdata                   (mm_interconnect_0_leds1_wr_val_s1_readdata),                  //                                     .readdata
		.leds1_wr_val_s1_writedata                  (mm_interconnect_0_leds1_wr_val_s1_writedata),                 //                                     .writedata
		.leds1_wr_val_s1_chipselect                 (mm_interconnect_0_leds1_wr_val_s1_chipselect),                //                                     .chipselect
		.leds2_brightness_s1_address                (mm_interconnect_0_leds2_brightness_s1_address),               //                  leds2_brightness_s1.address
		.leds2_brightness_s1_write                  (mm_interconnect_0_leds2_brightness_s1_write),                 //                                     .write
		.leds2_brightness_s1_readdata               (mm_interconnect_0_leds2_brightness_s1_readdata),              //                                     .readdata
		.leds2_brightness_s1_writedata              (mm_interconnect_0_leds2_brightness_s1_writedata),             //                                     .writedata
		.leds2_brightness_s1_chipselect             (mm_interconnect_0_leds2_brightness_s1_chipselect),            //                                     .chipselect
		.leds2_counter_s1_address                   (mm_interconnect_0_leds2_counter_s1_address),                  //                     leds2_counter_s1.address
		.leds2_counter_s1_readdata                  (mm_interconnect_0_leds2_counter_s1_readdata),                 //                                     .readdata
		.leds2_counter_of_s1_address                (mm_interconnect_0_leds2_counter_of_s1_address),               //                  leds2_counter_of_s1.address
		.leds2_counter_of_s1_readdata               (mm_interconnect_0_leds2_counter_of_s1_readdata),              //                                     .readdata
		.leds2_reset_control_s1_address             (mm_interconnect_0_leds2_reset_control_s1_address),            //               leds2_reset_control_s1.address
		.leds2_reset_control_s1_write               (mm_interconnect_0_leds2_reset_control_s1_write),              //                                     .write
		.leds2_reset_control_s1_readdata            (mm_interconnect_0_leds2_reset_control_s1_readdata),           //                                     .readdata
		.leds2_reset_control_s1_writedata           (mm_interconnect_0_leds2_reset_control_s1_writedata),          //                                     .writedata
		.leds2_reset_control_s1_chipselect          (mm_interconnect_0_leds2_reset_control_s1_chipselect),         //                                     .chipselect
		.leds2_wr_val_s1_address                    (mm_interconnect_0_leds2_wr_val_s1_address),                   //                      leds2_wr_val_s1.address
		.leds2_wr_val_s1_write                      (mm_interconnect_0_leds2_wr_val_s1_write),                     //                                     .write
		.leds2_wr_val_s1_readdata                   (mm_interconnect_0_leds2_wr_val_s1_readdata),                  //                                     .readdata
		.leds2_wr_val_s1_writedata                  (mm_interconnect_0_leds2_wr_val_s1_writedata),                 //                                     .writedata
		.leds2_wr_val_s1_chipselect                 (mm_interconnect_0_leds2_wr_val_s1_chipselect),                //                                     .chipselect
		.nios2e_jtag_debug_module_address           (mm_interconnect_0_nios2e_jtag_debug_module_address),          //             nios2e_jtag_debug_module.address
		.nios2e_jtag_debug_module_write             (mm_interconnect_0_nios2e_jtag_debug_module_write),            //                                     .write
		.nios2e_jtag_debug_module_read              (mm_interconnect_0_nios2e_jtag_debug_module_read),             //                                     .read
		.nios2e_jtag_debug_module_readdata          (mm_interconnect_0_nios2e_jtag_debug_module_readdata),         //                                     .readdata
		.nios2e_jtag_debug_module_writedata         (mm_interconnect_0_nios2e_jtag_debug_module_writedata),        //                                     .writedata
		.nios2e_jtag_debug_module_byteenable        (mm_interconnect_0_nios2e_jtag_debug_module_byteenable),       //                                     .byteenable
		.nios2e_jtag_debug_module_waitrequest       (mm_interconnect_0_nios2e_jtag_debug_module_waitrequest),      //                                     .waitrequest
		.nios2e_jtag_debug_module_debugaccess       (mm_interconnect_0_nios2e_jtag_debug_module_debugaccess),      //                                     .debugaccess
		.onchip_ram_s1_address                      (mm_interconnect_0_onchip_ram_s1_address),                     //                        onchip_ram_s1.address
		.onchip_ram_s1_write                        (mm_interconnect_0_onchip_ram_s1_write),                       //                                     .write
		.onchip_ram_s1_readdata                     (mm_interconnect_0_onchip_ram_s1_readdata),                    //                                     .readdata
		.onchip_ram_s1_writedata                    (mm_interconnect_0_onchip_ram_s1_writedata),                   //                                     .writedata
		.onchip_ram_s1_byteenable                   (mm_interconnect_0_onchip_ram_s1_byteenable),                  //                                     .byteenable
		.onchip_ram_s1_chipselect                   (mm_interconnect_0_onchip_ram_s1_chipselect),                  //                                     .chipselect
		.onchip_ram_s1_clken                        (mm_interconnect_0_onchip_ram_s1_clken),                       //                                     .clken
		.rc1_control_s1_address                     (mm_interconnect_0_rc1_control_s1_address),                    //                       rc1_control_s1.address
		.rc1_control_s1_write                       (mm_interconnect_0_rc1_control_s1_write),                      //                                     .write
		.rc1_control_s1_readdata                    (mm_interconnect_0_rc1_control_s1_readdata),                   //                                     .readdata
		.rc1_control_s1_writedata                   (mm_interconnect_0_rc1_control_s1_writedata),                  //                                     .writedata
		.rc1_control_s1_chipselect                  (mm_interconnect_0_rc1_control_s1_chipselect),                 //                                     .chipselect
		.rc1_ready_s1_address                       (mm_interconnect_0_rc1_ready_s1_address),                      //                         rc1_ready_s1.address
		.rc1_ready_s1_write                         (mm_interconnect_0_rc1_ready_s1_write),                        //                                     .write
		.rc1_ready_s1_readdata                      (mm_interconnect_0_rc1_ready_s1_readdata),                     //                                     .readdata
		.rc1_ready_s1_writedata                     (mm_interconnect_0_rc1_ready_s1_writedata),                    //                                     .writedata
		.rc1_ready_s1_chipselect                    (mm_interconnect_0_rc1_ready_s1_chipselect),                   //                                     .chipselect
		.sseg_brightness_s1_address                 (mm_interconnect_0_sseg_brightness_s1_address),                //                   sseg_brightness_s1.address
		.sseg_brightness_s1_write                   (mm_interconnect_0_sseg_brightness_s1_write),                  //                                     .write
		.sseg_brightness_s1_readdata                (mm_interconnect_0_sseg_brightness_s1_readdata),               //                                     .readdata
		.sseg_brightness_s1_writedata               (mm_interconnect_0_sseg_brightness_s1_writedata),              //                                     .writedata
		.sseg_brightness_s1_chipselect              (mm_interconnect_0_sseg_brightness_s1_chipselect),             //                                     .chipselect
		.sseg_counter_s1_address                    (mm_interconnect_0_sseg_counter_s1_address),                   //                      sseg_counter_s1.address
		.sseg_counter_s1_readdata                   (mm_interconnect_0_sseg_counter_s1_readdata),                  //                                     .readdata
		.sseg_counter_of_s1_address                 (mm_interconnect_0_sseg_counter_of_s1_address),                //                   sseg_counter_of_s1.address
		.sseg_counter_of_s1_readdata                (mm_interconnect_0_sseg_counter_of_s1_readdata),               //                                     .readdata
		.sseg_reset_control_s1_address              (mm_interconnect_0_sseg_reset_control_s1_address),             //                sseg_reset_control_s1.address
		.sseg_reset_control_s1_write                (mm_interconnect_0_sseg_reset_control_s1_write),               //                                     .write
		.sseg_reset_control_s1_readdata             (mm_interconnect_0_sseg_reset_control_s1_readdata),            //                                     .readdata
		.sseg_reset_control_s1_writedata            (mm_interconnect_0_sseg_reset_control_s1_writedata),           //                                     .writedata
		.sseg_reset_control_s1_chipselect           (mm_interconnect_0_sseg_reset_control_s1_chipselect),          //                                     .chipselect
		.sseg_wr_val_s1_address                     (mm_interconnect_0_sseg_wr_val_s1_address),                    //                       sseg_wr_val_s1.address
		.sseg_wr_val_s1_write                       (mm_interconnect_0_sseg_wr_val_s1_write),                      //                                     .write
		.sseg_wr_val_s1_readdata                    (mm_interconnect_0_sseg_wr_val_s1_readdata),                   //                                     .readdata
		.sseg_wr_val_s1_writedata                   (mm_interconnect_0_sseg_wr_val_s1_writedata),                  //                                     .writedata
		.sseg_wr_val_s1_chipselect                  (mm_interconnect_0_sseg_wr_val_s1_chipselect),                 //                                     .chipselect
		.status_led_en_s1_address                   (mm_interconnect_0_status_led_en_s1_address),                  //                     status_led_en_s1.address
		.status_led_en_s1_write                     (mm_interconnect_0_status_led_en_s1_write),                    //                                     .write
		.status_led_en_s1_readdata                  (mm_interconnect_0_status_led_en_s1_readdata),                 //                                     .readdata
		.status_led_en_s1_writedata                 (mm_interconnect_0_status_led_en_s1_writedata),                //                                     .writedata
		.status_led_en_s1_chipselect                (mm_interconnect_0_status_led_en_s1_chipselect),               //                                     .chipselect
		.sysid_c001_control_slave_address           (mm_interconnect_0_sysid_c001_control_slave_address),          //             sysid_c001_control_slave.address
		.sysid_c001_control_slave_readdata          (mm_interconnect_0_sysid_c001_control_slave_readdata),         //                                     .readdata
		.tc1_m_s1_address                           (mm_interconnect_0_tc1_m_s1_address),                          //                             tc1_m_s1.address
		.tc1_m_s1_write                             (mm_interconnect_0_tc1_m_s1_write),                            //                                     .write
		.tc1_m_s1_readdata                          (mm_interconnect_0_tc1_m_s1_readdata),                         //                                     .readdata
		.tc1_m_s1_writedata                         (mm_interconnect_0_tc1_m_s1_writedata),                        //                                     .writedata
		.tc1_m_s1_chipselect                        (mm_interconnect_0_tc1_m_s1_chipselect),                       //                                     .chipselect
		.tc1_status_s1_address                      (mm_interconnect_0_tc1_status_s1_address),                     //                        tc1_status_s1.address
		.tc1_status_s1_readdata                     (mm_interconnect_0_tc1_status_s1_readdata),                    //                                     .readdata
		.tc2_m_s1_address                           (mm_interconnect_0_tc2_m_s1_address),                          //                             tc2_m_s1.address
		.tc2_m_s1_write                             (mm_interconnect_0_tc2_m_s1_write),                            //                                     .write
		.tc2_m_s1_readdata                          (mm_interconnect_0_tc2_m_s1_readdata),                         //                                     .readdata
		.tc2_m_s1_writedata                         (mm_interconnect_0_tc2_m_s1_writedata),                        //                                     .writedata
		.tc2_m_s1_chipselect                        (mm_interconnect_0_tc2_m_s1_chipselect),                       //                                     .chipselect
		.tc2_status_s1_address                      (mm_interconnect_0_tc2_status_s1_address),                     //                        tc2_status_s1.address
		.tc2_status_s1_readdata                     (mm_interconnect_0_tc2_status_s1_readdata),                    //                                     .readdata
		.tc3_m_s1_address                           (mm_interconnect_0_tc3_m_s1_address),                          //                             tc3_m_s1.address
		.tc3_m_s1_write                             (mm_interconnect_0_tc3_m_s1_write),                            //                                     .write
		.tc3_m_s1_readdata                          (mm_interconnect_0_tc3_m_s1_readdata),                         //                                     .readdata
		.tc3_m_s1_writedata                         (mm_interconnect_0_tc3_m_s1_writedata),                        //                                     .writedata
		.tc3_m_s1_chipselect                        (mm_interconnect_0_tc3_m_s1_chipselect),                       //                                     .chipselect
		.tc3_status_s1_address                      (mm_interconnect_0_tc3_status_s1_address),                     //                        tc3_status_s1.address
		.tc3_status_s1_readdata                     (mm_interconnect_0_tc3_status_s1_readdata),                    //                                     .readdata
		.tc4_m_s1_address                           (mm_interconnect_0_tc4_m_s1_address),                          //                             tc4_m_s1.address
		.tc4_m_s1_write                             (mm_interconnect_0_tc4_m_s1_write),                            //                                     .write
		.tc4_m_s1_readdata                          (mm_interconnect_0_tc4_m_s1_readdata),                         //                                     .readdata
		.tc4_m_s1_writedata                         (mm_interconnect_0_tc4_m_s1_writedata),                        //                                     .writedata
		.tc4_m_s1_chipselect                        (mm_interconnect_0_tc4_m_s1_chipselect),                       //                                     .chipselect
		.tc4_status_s1_address                      (mm_interconnect_0_tc4_status_s1_address),                     //                        tc4_status_s1.address
		.tc4_status_s1_readdata                     (mm_interconnect_0_tc4_status_s1_readdata),                    //                                     .readdata
		.tc_reset_control_s1_address                (mm_interconnect_0_tc_reset_control_s1_address),               //                  tc_reset_control_s1.address
		.tc_reset_control_s1_write                  (mm_interconnect_0_tc_reset_control_s1_write),                 //                                     .write
		.tc_reset_control_s1_readdata               (mm_interconnect_0_tc_reset_control_s1_readdata),              //                                     .readdata
		.tc_reset_control_s1_writedata              (mm_interconnect_0_tc_reset_control_s1_writedata),             //                                     .writedata
		.tc_reset_control_s1_chipselect             (mm_interconnect_0_tc_reset_control_s1_chipselect),            //                                     .chipselect
		.uart1_baud_control_s1_address              (mm_interconnect_0_uart1_baud_control_s1_address),             //                uart1_baud_control_s1.address
		.uart1_baud_control_s1_write                (mm_interconnect_0_uart1_baud_control_s1_write),               //                                     .write
		.uart1_baud_control_s1_readdata             (mm_interconnect_0_uart1_baud_control_s1_readdata),            //                                     .readdata
		.uart1_baud_control_s1_writedata            (mm_interconnect_0_uart1_baud_control_s1_writedata),           //                                     .writedata
		.uart1_baud_control_s1_chipselect           (mm_interconnect_0_uart1_baud_control_s1_chipselect),          //                                     .chipselect
		.uart1_dvsr_s1_address                      (mm_interconnect_0_uart1_dvsr_s1_address),                     //                        uart1_dvsr_s1.address
		.uart1_dvsr_s1_write                        (mm_interconnect_0_uart1_dvsr_s1_write),                       //                                     .write
		.uart1_dvsr_s1_readdata                     (mm_interconnect_0_uart1_dvsr_s1_readdata),                    //                                     .readdata
		.uart1_dvsr_s1_writedata                    (mm_interconnect_0_uart1_dvsr_s1_writedata),                   //                                     .writedata
		.uart1_dvsr_s1_chipselect                   (mm_interconnect_0_uart1_dvsr_s1_chipselect),                  //                                     .chipselect
		.uart1_r_data_s1_address                    (mm_interconnect_0_uart1_r_data_s1_address),                   //                      uart1_r_data_s1.address
		.uart1_r_data_s1_readdata                   (mm_interconnect_0_uart1_r_data_s1_readdata),                  //                                     .readdata
		.uart1_reset_control_s1_address             (mm_interconnect_0_uart1_reset_control_s1_address),            //               uart1_reset_control_s1.address
		.uart1_reset_control_s1_write               (mm_interconnect_0_uart1_reset_control_s1_write),              //                                     .write
		.uart1_reset_control_s1_readdata            (mm_interconnect_0_uart1_reset_control_s1_readdata),           //                                     .readdata
		.uart1_reset_control_s1_writedata           (mm_interconnect_0_uart1_reset_control_s1_writedata),          //                                     .writedata
		.uart1_reset_control_s1_chipselect          (mm_interconnect_0_uart1_reset_control_s1_chipselect),         //                                     .chipselect
		.uart1_rx_counter_s1_address                (mm_interconnect_0_uart1_rx_counter_s1_address),               //                  uart1_rx_counter_s1.address
		.uart1_rx_counter_s1_readdata               (mm_interconnect_0_uart1_rx_counter_s1_readdata),              //                                     .readdata
		.uart1_status_control_s1_address            (mm_interconnect_0_uart1_status_control_s1_address),           //              uart1_status_control_s1.address
		.uart1_status_control_s1_readdata           (mm_interconnect_0_uart1_status_control_s1_readdata),          //                                     .readdata
		.uart1_tx_counter_s1_address                (mm_interconnect_0_uart1_tx_counter_s1_address),               //                  uart1_tx_counter_s1.address
		.uart1_tx_counter_s1_readdata               (mm_interconnect_0_uart1_tx_counter_s1_readdata),              //                                     .readdata
		.uart1_w_data_s1_address                    (mm_interconnect_0_uart1_w_data_s1_address),                   //                      uart1_w_data_s1.address
		.uart1_w_data_s1_write                      (mm_interconnect_0_uart1_w_data_s1_write),                     //                                     .write
		.uart1_w_data_s1_readdata                   (mm_interconnect_0_uart1_w_data_s1_readdata),                  //                                     .readdata
		.uart1_w_data_s1_writedata                  (mm_interconnect_0_uart1_w_data_s1_writedata),                 //                                     .writedata
		.uart1_w_data_s1_chipselect                 (mm_interconnect_0_uart1_w_data_s1_chipselect),                //                                     .chipselect
		.uart1_wr_control_s1_address                (mm_interconnect_0_uart1_wr_control_s1_address),               //                  uart1_wr_control_s1.address
		.uart1_wr_control_s1_write                  (mm_interconnect_0_uart1_wr_control_s1_write),                 //                                     .write
		.uart1_wr_control_s1_readdata               (mm_interconnect_0_uart1_wr_control_s1_readdata),              //                                     .readdata
		.uart1_wr_control_s1_writedata              (mm_interconnect_0_uart1_wr_control_s1_writedata),             //                                     .writedata
		.uart1_wr_control_s1_chipselect             (mm_interconnect_0_uart1_wr_control_s1_chipselect),            //                                     .chipselect
		.warn_pwm_brightness_s1_address             (mm_interconnect_0_warn_pwm_brightness_s1_address),            //               warn_pwm_brightness_s1.address
		.warn_pwm_brightness_s1_write               (mm_interconnect_0_warn_pwm_brightness_s1_write),              //                                     .write
		.warn_pwm_brightness_s1_readdata            (mm_interconnect_0_warn_pwm_brightness_s1_readdata),           //                                     .readdata
		.warn_pwm_brightness_s1_writedata           (mm_interconnect_0_warn_pwm_brightness_s1_writedata),          //                                     .writedata
		.warn_pwm_brightness_s1_chipselect          (mm_interconnect_0_warn_pwm_brightness_s1_chipselect),         //                                     .chipselect
		.warn_pwm_control_s1_address                (mm_interconnect_0_warn_pwm_control_s1_address),               //                  warn_pwm_control_s1.address
		.warn_pwm_control_s1_write                  (mm_interconnect_0_warn_pwm_control_s1_write),                 //                                     .write
		.warn_pwm_control_s1_readdata               (mm_interconnect_0_warn_pwm_control_s1_readdata),              //                                     .readdata
		.warn_pwm_control_s1_writedata              (mm_interconnect_0_warn_pwm_control_s1_writedata),             //                                     .writedata
		.warn_pwm_control_s1_chipselect             (mm_interconnect_0_warn_pwm_control_s1_chipselect)             //                                     .chipselect
	);

	controller_irq_mapper irq_mapper (
		.clk           (clock_50_clk),                   //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (nios2e_d_irq_irq)                //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                       // reset_in0.reset
		.reset_in1      (nios2e_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clock_50_clk),                         //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),       // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),   //          .reset_req
		.reset_req_in0  (1'b0),                                 // (terminated)
		.reset_req_in1  (1'b0),                                 // (terminated)
		.reset_in2      (1'b0),                                 // (terminated)
		.reset_req_in2  (1'b0),                                 // (terminated)
		.reset_in3      (1'b0),                                 // (terminated)
		.reset_req_in3  (1'b0),                                 // (terminated)
		.reset_in4      (1'b0),                                 // (terminated)
		.reset_req_in4  (1'b0),                                 // (terminated)
		.reset_in5      (1'b0),                                 // (terminated)
		.reset_req_in5  (1'b0),                                 // (terminated)
		.reset_in6      (1'b0),                                 // (terminated)
		.reset_req_in6  (1'b0),                                 // (terminated)
		.reset_in7      (1'b0),                                 // (terminated)
		.reset_req_in7  (1'b0),                                 // (terminated)
		.reset_in8      (1'b0),                                 // (terminated)
		.reset_req_in8  (1'b0),                                 // (terminated)
		.reset_in9      (1'b0),                                 // (terminated)
		.reset_req_in9  (1'b0),                                 // (terminated)
		.reset_in10     (1'b0),                                 // (terminated)
		.reset_req_in10 (1'b0),                                 // (terminated)
		.reset_in11     (1'b0),                                 // (terminated)
		.reset_req_in11 (1'b0),                                 // (terminated)
		.reset_in12     (1'b0),                                 // (terminated)
		.reset_req_in12 (1'b0),                                 // (terminated)
		.reset_in13     (1'b0),                                 // (terminated)
		.reset_req_in13 (1'b0),                                 // (terminated)
		.reset_in14     (1'b0),                                 // (terminated)
		.reset_req_in14 (1'b0),                                 // (terminated)
		.reset_in15     (1'b0),                                 // (terminated)
		.reset_req_in15 (1'b0)                                  // (terminated)
	);

endmodule
